module u_cla(input [7:0] a, input [7:0] b, output [8:0] u_cla_out);
  wire u_cla_pg_logic0_pg_logic_or0;
  wire u_cla_pg_logic0_pg_logic_and0;
  wire u_cla_pg_logic0_pg_logic_xor0;
  wire u_cla_pg_logic1_pg_logic_or0;
  wire u_cla_pg_logic1_pg_logic_and0;
  wire u_cla_pg_logic1_pg_logic_xor0;
  wire u_cla_xor1;
  wire u_cla_and0_1_1_0_0;
  wire u_cla_or0_1_1_0;
  wire u_cla_pg_logic2_pg_logic_or0;
  wire u_cla_pg_logic2_pg_logic_and0;
  wire u_cla_pg_logic2_pg_logic_xor0;
  wire u_cla_xor2;
  wire u_cla_and0_2_0_1_1;
  wire u_cla_and0_2_1_0_2;
  wire u_cla_and0_2_1_1_3;
  wire u_cla_and0_2_2_0_4;
  wire u_cla_orred0_2_2__1_1;
  wire u_cla_or0_2_2_2;
  wire u_cla_pg_logic3_pg_logic_or0;
  wire u_cla_pg_logic3_pg_logic_and0;
  wire u_cla_pg_logic3_pg_logic_xor0;
  wire u_cla_xor3;
  wire u_cla_and0_3_0_1_5;
  wire u_cla_and0_3_1_0_6;
  wire u_cla_and0_3_1_1_7;
  wire u_cla_and0_3_1_2_8;
  wire u_cla_and0_3_2_0_9;
  wire u_cla_and0_3_2_1_10;
  wire u_cla_and0_3_3_0_11;
  wire u_cla_orred0_3_3__1_3;
  wire u_cla_orred0_3_3__2_4;
  wire u_cla_or0_3_3_5;
  wire u_cla_pg_logic4_pg_logic_or0;
  wire u_cla_pg_logic4_pg_logic_and0;
  wire u_cla_pg_logic4_pg_logic_xor0;
  wire u_cla_xor4;
  wire u_cla_and1_0_0_0_12;
  wire u_cla_or1_0_0_6;
  wire u_cla_pg_logic5_pg_logic_or0;
  wire u_cla_pg_logic5_pg_logic_and0;
  wire u_cla_pg_logic5_pg_logic_xor0;
  wire u_cla_xor5;
  wire u_cla_and1_1_0_0_13;
  wire u_cla_and1_1_0_1_14;
  wire u_cla_and1_1_1_0_15;
  wire u_cla_orred1_1_1__0_7;
  wire u_cla_or1_1_1_8;
  wire u_cla_pg_logic6_pg_logic_or0;
  wire u_cla_pg_logic6_pg_logic_and0;
  wire u_cla_pg_logic6_pg_logic_xor0;
  wire u_cla_xor6;
  wire u_cla_and1_2_0_0_16;
  wire u_cla_and1_2_0_1_17;
  wire u_cla_and1_2_0_2_18;
  wire u_cla_and1_2_1_0_19;
  wire u_cla_and1_2_1_1_20;
  wire u_cla_and1_2_2_0_21;
  wire u_cla_orred1_2_2__0_9;
  wire u_cla_orred1_2_2__1_10;
  wire u_cla_or1_2_2_11;
  wire u_cla_pg_logic7_pg_logic_or0;
  wire u_cla_pg_logic7_pg_logic_and0;
  wire u_cla_pg_logic7_pg_logic_xor0;
  wire u_cla_xor7;
  wire u_cla_and1_3_0_0_22;
  wire u_cla_and1_3_0_1_23;
  wire u_cla_and1_3_0_2_24;
  wire u_cla_and1_3_0_3_25;
  wire u_cla_and1_3_1_0_26;
  wire u_cla_and1_3_1_1_27;
  wire u_cla_and1_3_1_2_28;
  wire u_cla_and1_3_2_0_29;
  wire u_cla_and1_3_2_1_30;
  wire u_cla_and1_3_3_0_31;
  wire u_cla_orred1_3_3__0_12;
  wire u_cla_orred1_3_3__1_13;
  wire u_cla_orred1_3_3__2_14;
  wire u_cla_or1_3_3_15;

  assign u_cla_pg_logic0_pg_logic_or0 = a[0] | b[0];
  assign u_cla_pg_logic0_pg_logic_and0 = a[0] & b[0];
  assign u_cla_pg_logic0_pg_logic_xor0 = a[0] ^ b[0];
  assign u_cla_pg_logic1_pg_logic_or0 = a[1] | b[1];
  assign u_cla_pg_logic1_pg_logic_and0 = a[1] & b[1];
  assign u_cla_pg_logic1_pg_logic_xor0 = a[1] ^ b[1];
  assign u_cla_xor1 = u_cla_pg_logic1_pg_logic_xor0 ^ u_cla_pg_logic0_pg_logic_and0;
  assign u_cla_and0_1_1_0_0 = u_cla_pg_logic0_pg_logic_and0 & u_cla_pg_logic1_pg_logic_or0;
  assign u_cla_or0_1_1_0 = u_cla_pg_logic1_pg_logic_and0 | u_cla_and0_1_1_0_0;
  assign u_cla_pg_logic2_pg_logic_or0 = a[2] | b[2];
  assign u_cla_pg_logic2_pg_logic_and0 = a[2] & b[2];
  assign u_cla_pg_logic2_pg_logic_xor0 = a[2] ^ b[2];
  assign u_cla_xor2 = u_cla_pg_logic2_pg_logic_xor0 ^ u_cla_or0_1_1_0;
  assign u_cla_and0_2_0_1_1 = u_cla_pg_logic2_pg_logic_or0 & u_cla_pg_logic0_pg_logic_or0;
  assign u_cla_and0_2_1_0_2 = u_cla_pg_logic0_pg_logic_and0 & u_cla_pg_logic2_pg_logic_or0;
  assign u_cla_and0_2_1_1_3 = u_cla_and0_2_1_0_2 & u_cla_pg_logic1_pg_logic_or0;
  assign u_cla_and0_2_2_0_4 = u_cla_pg_logic1_pg_logic_and0 & u_cla_pg_logic2_pg_logic_or0;
  assign u_cla_orred0_2_2__1_1 = u_cla_and0_2_1_1_3 | u_cla_and0_2_2_0_4;
  assign u_cla_or0_2_2_2 = u_cla_pg_logic2_pg_logic_and0 | u_cla_orred0_2_2__1_1;
  assign u_cla_pg_logic3_pg_logic_or0 = a[3] | b[3];
  assign u_cla_pg_logic3_pg_logic_and0 = a[3] & b[3];
  assign u_cla_pg_logic3_pg_logic_xor0 = a[3] ^ b[3];
  assign u_cla_xor3 = u_cla_pg_logic3_pg_logic_xor0 ^ u_cla_or0_2_2_2;
  assign u_cla_and0_3_0_1_5 = u_cla_pg_logic3_pg_logic_or0 & u_cla_pg_logic1_pg_logic_or0;
  assign u_cla_and0_3_1_0_6 = u_cla_pg_logic0_pg_logic_and0 & u_cla_pg_logic2_pg_logic_or0;
  assign u_cla_and0_3_1_1_7 = u_cla_pg_logic3_pg_logic_or0 & u_cla_pg_logic1_pg_logic_or0;
  assign u_cla_and0_3_1_2_8 = u_cla_and0_3_1_0_6 & u_cla_and0_3_1_1_7;
  assign u_cla_and0_3_2_0_9 = u_cla_pg_logic1_pg_logic_and0 & u_cla_pg_logic3_pg_logic_or0;
  assign u_cla_and0_3_2_1_10 = u_cla_and0_3_2_0_9 & u_cla_pg_logic2_pg_logic_or0;
  assign u_cla_and0_3_3_0_11 = u_cla_pg_logic2_pg_logic_and0 & u_cla_pg_logic3_pg_logic_or0;
  assign u_cla_orred0_3_3__1_3 = u_cla_and0_3_1_2_8 | u_cla_and0_3_3_0_11;
  assign u_cla_orred0_3_3__2_4 = u_cla_and0_3_2_1_10 | u_cla_orred0_3_3__1_3;
  assign u_cla_or0_3_3_5 = u_cla_pg_logic3_pg_logic_and0 | u_cla_orred0_3_3__2_4;
  assign u_cla_pg_logic4_pg_logic_or0 = a[4] | b[4];
  assign u_cla_pg_logic4_pg_logic_and0 = a[4] & b[4];
  assign u_cla_pg_logic4_pg_logic_xor0 = a[4] ^ b[4];
  assign u_cla_xor4 = u_cla_pg_logic4_pg_logic_xor0 ^ u_cla_or0_3_3_5;
  assign u_cla_and1_0_0_0_12 = u_cla_or0_3_3_5 & u_cla_pg_logic4_pg_logic_or0;
  assign u_cla_or1_0_0_6 = u_cla_pg_logic4_pg_logic_and0 | u_cla_and1_0_0_0_12;
  assign u_cla_pg_logic5_pg_logic_or0 = a[5] | b[5];
  assign u_cla_pg_logic5_pg_logic_and0 = a[5] & b[5];
  assign u_cla_pg_logic5_pg_logic_xor0 = a[5] ^ b[5];
  assign u_cla_xor5 = u_cla_pg_logic5_pg_logic_xor0 ^ u_cla_or1_0_0_6;
  assign u_cla_and1_1_0_0_13 = u_cla_or0_3_3_5 & u_cla_pg_logic5_pg_logic_or0;
  assign u_cla_and1_1_0_1_14 = u_cla_and1_1_0_0_13 & u_cla_pg_logic4_pg_logic_or0;
  assign u_cla_and1_1_1_0_15 = u_cla_pg_logic4_pg_logic_and0 & u_cla_pg_logic5_pg_logic_or0;
  assign u_cla_orred1_1_1__0_7 = u_cla_and1_1_0_1_14 | u_cla_and1_1_1_0_15;
  assign u_cla_or1_1_1_8 = u_cla_pg_logic5_pg_logic_and0 | u_cla_orred1_1_1__0_7;
  assign u_cla_pg_logic6_pg_logic_or0 = a[6] | b[6];
  assign u_cla_pg_logic6_pg_logic_and0 = a[6] & b[6];
  assign u_cla_pg_logic6_pg_logic_xor0 = a[6] ^ b[6];
  assign u_cla_xor6 = u_cla_pg_logic6_pg_logic_xor0 ^ u_cla_or1_1_1_8;
  assign u_cla_and1_2_0_0_16 = u_cla_or0_3_3_5 & u_cla_pg_logic5_pg_logic_or0;
  assign u_cla_and1_2_0_1_17 = u_cla_pg_logic6_pg_logic_or0 & u_cla_pg_logic4_pg_logic_or0;
  assign u_cla_and1_2_0_2_18 = u_cla_and1_2_0_0_16 & u_cla_and1_2_0_1_17;
  assign u_cla_and1_2_1_0_19 = u_cla_pg_logic4_pg_logic_and0 & u_cla_pg_logic6_pg_logic_or0;
  assign u_cla_and1_2_1_1_20 = u_cla_and1_2_1_0_19 & u_cla_pg_logic5_pg_logic_or0;
  assign u_cla_and1_2_2_0_21 = u_cla_pg_logic5_pg_logic_and0 & u_cla_pg_logic6_pg_logic_or0;
  assign u_cla_orred1_2_2__0_9 = u_cla_and1_2_0_2_18 | u_cla_and1_2_1_1_20;
  assign u_cla_orred1_2_2__1_10 = u_cla_orred1_2_2__0_9 | u_cla_and1_2_2_0_21;
  assign u_cla_or1_2_2_11 = u_cla_pg_logic6_pg_logic_and0 | u_cla_orred1_2_2__1_10;
  assign u_cla_pg_logic7_pg_logic_or0 = a[7] | b[7];
  assign u_cla_pg_logic7_pg_logic_and0 = a[7] & b[7];
  assign u_cla_pg_logic7_pg_logic_xor0 = a[7] ^ b[7];
  assign u_cla_xor7 = u_cla_pg_logic7_pg_logic_xor0 ^ u_cla_or1_2_2_11;
  assign u_cla_and1_3_0_0_22 = u_cla_or0_3_3_5 & u_cla_pg_logic6_pg_logic_or0;
  assign u_cla_and1_3_0_1_23 = u_cla_pg_logic7_pg_logic_or0 & u_cla_pg_logic5_pg_logic_or0;
  assign u_cla_and1_3_0_2_24 = u_cla_and1_3_0_0_22 & u_cla_and1_3_0_1_23;
  assign u_cla_and1_3_0_3_25 = u_cla_and1_3_0_2_24 & u_cla_pg_logic4_pg_logic_or0;
  assign u_cla_and1_3_1_0_26 = u_cla_pg_logic4_pg_logic_and0 & u_cla_pg_logic6_pg_logic_or0;
  assign u_cla_and1_3_1_1_27 = u_cla_pg_logic7_pg_logic_or0 & u_cla_pg_logic5_pg_logic_or0;
  assign u_cla_and1_3_1_2_28 = u_cla_and1_3_1_0_26 & u_cla_and1_3_1_1_27;
  assign u_cla_and1_3_2_0_29 = u_cla_pg_logic5_pg_logic_and0 & u_cla_pg_logic7_pg_logic_or0;
  assign u_cla_and1_3_2_1_30 = u_cla_and1_3_2_0_29 & u_cla_pg_logic6_pg_logic_or0;
  assign u_cla_and1_3_3_0_31 = u_cla_pg_logic6_pg_logic_and0 & u_cla_pg_logic7_pg_logic_or0;
  assign u_cla_orred1_3_3__0_12 = u_cla_and1_3_0_3_25 | u_cla_and1_3_2_1_30;
  assign u_cla_orred1_3_3__1_13 = u_cla_and1_3_1_2_28 | u_cla_and1_3_3_0_31;
  assign u_cla_orred1_3_3__2_14 = u_cla_orred1_3_3__0_12 | u_cla_orred1_3_3__1_13;
  assign u_cla_or1_3_3_15 = u_cla_pg_logic7_pg_logic_and0 | u_cla_orred1_3_3__2_14;

  assign u_cla_out[0] = u_cla_pg_logic0_pg_logic_xor0;
  assign u_cla_out[1] = u_cla_xor1;
  assign u_cla_out[2] = u_cla_xor2;
  assign u_cla_out[3] = u_cla_xor3;
  assign u_cla_out[4] = u_cla_xor4;
  assign u_cla_out[5] = u_cla_xor5;
  assign u_cla_out[6] = u_cla_xor6;
  assign u_cla_out[7] = u_cla_xor7;
  assign u_cla_out[8] = u_cla_or1_3_3_15;
endmodule