module u_rca(input [7:0] a, input [7:0] b, output [8:0] u_rca_out);
  wire u_rca_ha_ha_xor0;
  wire u_rca_ha_ha_and0;
  wire u_rca_fa1_fa_xor0;
  wire u_rca_fa1_fa_and0;
  wire u_rca_fa1_fa_xor1;
  wire u_rca_fa1_fa_and1;
  wire u_rca_fa1_fa_or0;
  wire u_rca_fa2_fa_xor0;
  wire u_rca_fa2_fa_and0;
  wire u_rca_fa2_fa_xor1;
  wire u_rca_fa2_fa_and1;
  wire u_rca_fa2_fa_or0;
  wire u_rca_fa3_fa_xor0;
  wire u_rca_fa3_fa_and0;
  wire u_rca_fa3_fa_xor1;
  wire u_rca_fa3_fa_and1;
  wire u_rca_fa3_fa_or0;
  wire u_rca_fa4_fa_xor0;
  wire u_rca_fa4_fa_and0;
  wire u_rca_fa4_fa_xor1;
  wire u_rca_fa4_fa_and1;
  wire u_rca_fa4_fa_or0;
  wire u_rca_fa5_fa_xor0;
  wire u_rca_fa5_fa_and0;
  wire u_rca_fa5_fa_xor1;
  wire u_rca_fa5_fa_and1;
  wire u_rca_fa5_fa_or0;
  wire u_rca_fa6_fa_xor0;
  wire u_rca_fa6_fa_and0;
  wire u_rca_fa6_fa_xor1;
  wire u_rca_fa6_fa_and1;
  wire u_rca_fa6_fa_or0;
  wire u_rca_fa7_fa_xor0;
  wire u_rca_fa7_fa_and0;
  wire u_rca_fa7_fa_xor1;
  wire u_rca_fa7_fa_and1;
  wire u_rca_fa7_fa_or0;

  assign u_rca_ha_ha_xor0 = a[0] ^ b[0];
  assign u_rca_ha_ha_and0 = a[0] & b[0];
  assign u_rca_fa1_fa_xor0 = a[1] ^ b[1];
  assign u_rca_fa1_fa_and0 = a[1] & b[1];
  assign u_rca_fa1_fa_xor1 = u_rca_fa1_fa_xor0 ^ u_rca_ha_ha_and0;
  assign u_rca_fa1_fa_and1 = u_rca_fa1_fa_xor0 & u_rca_ha_ha_and0;
  assign u_rca_fa1_fa_or0 = u_rca_fa1_fa_and0 | u_rca_fa1_fa_and1;
  assign u_rca_fa2_fa_xor0 = a[2] ^ b[2];
  assign u_rca_fa2_fa_and0 = a[2] & b[2];
  assign u_rca_fa2_fa_xor1 = u_rca_fa2_fa_xor0 ^ u_rca_fa1_fa_or0;
  assign u_rca_fa2_fa_and1 = u_rca_fa2_fa_xor0 & u_rca_fa1_fa_or0;
  assign u_rca_fa2_fa_or0 = u_rca_fa2_fa_and0 | u_rca_fa2_fa_and1;
  assign u_rca_fa3_fa_xor0 = a[3] ^ b[3];
  assign u_rca_fa3_fa_and0 = a[3] & b[3];
  assign u_rca_fa3_fa_xor1 = u_rca_fa3_fa_xor0 ^ u_rca_fa2_fa_or0;
  assign u_rca_fa3_fa_and1 = u_rca_fa3_fa_xor0 & u_rca_fa2_fa_or0;
  assign u_rca_fa3_fa_or0 = u_rca_fa3_fa_and0 | u_rca_fa3_fa_and1;
  assign u_rca_fa4_fa_xor0 = a[4] ^ b[4];
  assign u_rca_fa4_fa_and0 = a[4] & b[4];
  assign u_rca_fa4_fa_xor1 = u_rca_fa4_fa_xor0 ^ u_rca_fa3_fa_or0;
  assign u_rca_fa4_fa_and1 = u_rca_fa4_fa_xor0 & u_rca_fa3_fa_or0;
  assign u_rca_fa4_fa_or0 = u_rca_fa4_fa_and0 | u_rca_fa4_fa_and1;
  assign u_rca_fa5_fa_xor0 = a[5] ^ b[5];
  assign u_rca_fa5_fa_and0 = a[5] & b[5];
  assign u_rca_fa5_fa_xor1 = u_rca_fa5_fa_xor0 ^ u_rca_fa4_fa_or0;
  assign u_rca_fa5_fa_and1 = u_rca_fa5_fa_xor0 & u_rca_fa4_fa_or0;
  assign u_rca_fa5_fa_or0 = u_rca_fa5_fa_and0 | u_rca_fa5_fa_and1;
  assign u_rca_fa6_fa_xor0 = a[6] ^ b[6];
  assign u_rca_fa6_fa_and0 = a[6] & b[6];
  assign u_rca_fa6_fa_xor1 = u_rca_fa6_fa_xor0 ^ u_rca_fa5_fa_or0;
  assign u_rca_fa6_fa_and1 = u_rca_fa6_fa_xor0 & u_rca_fa5_fa_or0;
  assign u_rca_fa6_fa_or0 = u_rca_fa6_fa_and0 | u_rca_fa6_fa_and1;
  assign u_rca_fa7_fa_xor0 = a[7] ^ b[7];
  assign u_rca_fa7_fa_and0 = a[7] & b[7];
  assign u_rca_fa7_fa_xor1 = u_rca_fa7_fa_xor0 ^ u_rca_fa6_fa_or0;
  assign u_rca_fa7_fa_and1 = u_rca_fa7_fa_xor0 & u_rca_fa6_fa_or0;
  assign u_rca_fa7_fa_or0 = u_rca_fa7_fa_and0 | u_rca_fa7_fa_and1;

  assign u_rca_out[0] = u_rca_ha_ha_xor0;
  assign u_rca_out[1] = u_rca_fa1_fa_xor1;
  assign u_rca_out[2] = u_rca_fa2_fa_xor1;
  assign u_rca_out[3] = u_rca_fa3_fa_xor1;
  assign u_rca_out[4] = u_rca_fa4_fa_xor1;
  assign u_rca_out[5] = u_rca_fa5_fa_xor1;
  assign u_rca_out[6] = u_rca_fa6_fa_xor1;
  assign u_rca_out[7] = u_rca_fa7_fa_xor1;
  assign u_rca_out[8] = u_rca_fa7_fa_or0;
endmodule