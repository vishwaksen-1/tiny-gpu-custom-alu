module u_rcs(input [7:0] a, input [7:0] b, output [8:0] u_rcs_out);
  wire u_rcs_not0;
  wire u_rcs_ha_fa_xor0;
  wire u_rcs_ha_fa_and0;
  wire u_rcs_ha_fa_xor1_not;
  wire u_rcs_ha_fa_or0;
  wire u_rcs_not1;
  wire u_rcs_fa1_fa_xor0;
  wire u_rcs_fa1_fa_and0;
  wire u_rcs_fa1_fa_xor1;
  wire u_rcs_fa1_fa_and1;
  wire u_rcs_fa1_fa_or0;
  wire u_rcs_not2;
  wire u_rcs_fa2_fa_xor0;
  wire u_rcs_fa2_fa_and0;
  wire u_rcs_fa2_fa_xor1;
  wire u_rcs_fa2_fa_and1;
  wire u_rcs_fa2_fa_or0;
  wire u_rcs_not3;
  wire u_rcs_fa3_fa_xor0;
  wire u_rcs_fa3_fa_and0;
  wire u_rcs_fa3_fa_xor1;
  wire u_rcs_fa3_fa_and1;
  wire u_rcs_fa3_fa_or0;
  wire u_rcs_not4;
  wire u_rcs_fa4_fa_xor0;
  wire u_rcs_fa4_fa_and0;
  wire u_rcs_fa4_fa_xor1;
  wire u_rcs_fa4_fa_and1;
  wire u_rcs_fa4_fa_or0;
  wire u_rcs_not5;
  wire u_rcs_fa5_fa_xor0;
  wire u_rcs_fa5_fa_and0;
  wire u_rcs_fa5_fa_xor1;
  wire u_rcs_fa5_fa_and1;
  wire u_rcs_fa5_fa_or0;
  wire u_rcs_not6;
  wire u_rcs_fa6_fa_xor0;
  wire u_rcs_fa6_fa_and0;
  wire u_rcs_fa6_fa_xor1;
  wire u_rcs_fa6_fa_and1;
  wire u_rcs_fa6_fa_or0;
  wire u_rcs_not7;
  wire u_rcs_fa7_fa_xor0;
  wire u_rcs_fa7_fa_and0;
  wire u_rcs_fa7_fa_xor1;
  wire u_rcs_fa7_fa_and1;
  wire u_rcs_fa7_fa_or0;
  wire u_rcs_not_c7;

  assign u_rcs_not0 = ~b[0];
  assign u_rcs_ha_fa_xor0 = a[0] ^ u_rcs_not0;
  assign u_rcs_ha_fa_and0 = a[0] & u_rcs_not0;
  assign u_rcs_ha_fa_xor1_not = ~u_rcs_ha_fa_xor0;
  assign u_rcs_ha_fa_or0 = u_rcs_ha_fa_and0 | u_rcs_ha_fa_xor0;
  assign u_rcs_not1 = ~b[1];
  assign u_rcs_fa1_fa_xor0 = a[1] ^ u_rcs_not1;
  assign u_rcs_fa1_fa_and0 = a[1] & u_rcs_not1;
  assign u_rcs_fa1_fa_xor1 = u_rcs_fa1_fa_xor0 ^ u_rcs_ha_fa_or0;
  assign u_rcs_fa1_fa_and1 = u_rcs_fa1_fa_xor0 & u_rcs_ha_fa_or0;
  assign u_rcs_fa1_fa_or0 = u_rcs_fa1_fa_and0 | u_rcs_fa1_fa_and1;
  assign u_rcs_not2 = ~b[2];
  assign u_rcs_fa2_fa_xor0 = a[2] ^ u_rcs_not2;
  assign u_rcs_fa2_fa_and0 = a[2] & u_rcs_not2;
  assign u_rcs_fa2_fa_xor1 = u_rcs_fa2_fa_xor0 ^ u_rcs_fa1_fa_or0;
  assign u_rcs_fa2_fa_and1 = u_rcs_fa2_fa_xor0 & u_rcs_fa1_fa_or0;
  assign u_rcs_fa2_fa_or0 = u_rcs_fa2_fa_and0 | u_rcs_fa2_fa_and1;
  assign u_rcs_not3 = ~b[3];
  assign u_rcs_fa3_fa_xor0 = a[3] ^ u_rcs_not3;
  assign u_rcs_fa3_fa_and0 = a[3] & u_rcs_not3;
  assign u_rcs_fa3_fa_xor1 = u_rcs_fa3_fa_xor0 ^ u_rcs_fa2_fa_or0;
  assign u_rcs_fa3_fa_and1 = u_rcs_fa3_fa_xor0 & u_rcs_fa2_fa_or0;
  assign u_rcs_fa3_fa_or0 = u_rcs_fa3_fa_and0 | u_rcs_fa3_fa_and1;
  assign u_rcs_not4 = ~b[4];
  assign u_rcs_fa4_fa_xor0 = a[4] ^ u_rcs_not4;
  assign u_rcs_fa4_fa_and0 = a[4] & u_rcs_not4;
  assign u_rcs_fa4_fa_xor1 = u_rcs_fa4_fa_xor0 ^ u_rcs_fa3_fa_or0;
  assign u_rcs_fa4_fa_and1 = u_rcs_fa4_fa_xor0 & u_rcs_fa3_fa_or0;
  assign u_rcs_fa4_fa_or0 = u_rcs_fa4_fa_and0 | u_rcs_fa4_fa_and1;
  assign u_rcs_not5 = ~b[5];
  assign u_rcs_fa5_fa_xor0 = a[5] ^ u_rcs_not5;
  assign u_rcs_fa5_fa_and0 = a[5] & u_rcs_not5;
  assign u_rcs_fa5_fa_xor1 = u_rcs_fa5_fa_xor0 ^ u_rcs_fa4_fa_or0;
  assign u_rcs_fa5_fa_and1 = u_rcs_fa5_fa_xor0 & u_rcs_fa4_fa_or0;
  assign u_rcs_fa5_fa_or0 = u_rcs_fa5_fa_and0 | u_rcs_fa5_fa_and1;
  assign u_rcs_not6 = ~b[6];
  assign u_rcs_fa6_fa_xor0 = a[6] ^ u_rcs_not6;
  assign u_rcs_fa6_fa_and0 = a[6] & u_rcs_not6;
  assign u_rcs_fa6_fa_xor1 = u_rcs_fa6_fa_xor0 ^ u_rcs_fa5_fa_or0;
  assign u_rcs_fa6_fa_and1 = u_rcs_fa6_fa_xor0 & u_rcs_fa5_fa_or0;
  assign u_rcs_fa6_fa_or0 = u_rcs_fa6_fa_and0 | u_rcs_fa6_fa_and1;
  assign u_rcs_not7 = ~b[7];
  assign u_rcs_fa7_fa_xor0 = a[7] ^ u_rcs_not7;
  assign u_rcs_fa7_fa_and0 = a[7] & u_rcs_not7;
  assign u_rcs_fa7_fa_xor1 = u_rcs_fa7_fa_xor0 ^ u_rcs_fa6_fa_or0;
  assign u_rcs_fa7_fa_and1 = u_rcs_fa7_fa_xor0 & u_rcs_fa6_fa_or0;
  assign u_rcs_fa7_fa_or0 = u_rcs_fa7_fa_and0 | u_rcs_fa7_fa_and1;
  assign u_rcs_not_c7 = ~u_rcs_fa7_fa_or0;

  assign u_rcs_out[0] = u_rcs_ha_fa_xor1_not;
  assign u_rcs_out[1] = u_rcs_fa1_fa_xor1;
  assign u_rcs_out[2] = u_rcs_fa2_fa_xor1;
  assign u_rcs_out[3] = u_rcs_fa3_fa_xor1;
  assign u_rcs_out[4] = u_rcs_fa4_fa_xor1;
  assign u_rcs_out[5] = u_rcs_fa5_fa_xor1;
  assign u_rcs_out[6] = u_rcs_fa6_fa_xor1;
  assign u_rcs_out[7] = u_rcs_fa7_fa_xor1;
  assign u_rcs_out[8] = u_rcs_not_c7;
endmodule