module u_cosa(input [7:0] a, input [7:0] b, output [8:0] u_cosa_out);
  wire u_cosa_fa0_fa_xor0;
  wire u_cosa_fa0_fa_and0;
  wire u_cosa_fa1_fa_xor0;
  wire u_cosa_fa1_fa_and0;
  wire u_cosa_fa2_fa_xor0;
  wire u_cosa_fa2_fa_and0;
  wire u_cosa_fa2_fa_xor1_not;
  wire u_cosa_fa2_fa_or0;
  wire u_cosa_mux2to1_0_mux2to1_and0;
  wire u_cosa_mux2to1_0_mux2to1_not0;
  wire u_cosa_mux2to1_0_mux2to1_and1;
  wire u_cosa_mux2to1_0_mux2to1_xor0;
  wire u_cosa_mux2to1_1_mux2to1_and0;
  wire u_cosa_mux2to1_1_mux2to1_not0;
  wire u_cosa_mux2to1_1_mux2to1_and1;
  wire u_cosa_mux2to1_1_mux2to1_xor0;
  wire u_cosa_fa3_fa_xor0;
  wire u_cosa_fa3_fa_and0;
  wire u_cosa_fa4_fa_xor0;
  wire u_cosa_fa4_fa_and0;
  wire u_cosa_fa4_fa_xor1_not;
  wire u_cosa_fa4_fa_or0;
  wire u_cosa_mux2to1_2_mux2to1_and0;
  wire u_cosa_mux2to1_2_mux2to1_not0;
  wire u_cosa_mux2to1_2_mux2to1_and1;
  wire u_cosa_mux2to1_2_mux2to1_xor0;
  wire u_cosa_fa5_fa_xor0;
  wire u_cosa_fa5_fa_and0;
  wire u_cosa_fa6_fa_xor0;
  wire u_cosa_fa6_fa_and0;
  wire u_cosa_fa6_fa_xor1_not;
  wire u_cosa_fa6_fa_or0;
  wire u_cosa_mux2to1_3_mux2to1_and0;
  wire u_cosa_mux2to1_3_mux2to1_not0;
  wire u_cosa_mux2to1_3_mux2to1_and1;
  wire u_cosa_mux2to1_3_mux2to1_xor0;
  wire u_cosa_mux2to1_4_mux2to1_and0;
  wire u_cosa_mux2to1_4_mux2to1_not0;
  wire u_cosa_mux2to1_4_mux2to1_and1;
  wire u_cosa_mux2to1_4_mux2to1_xor0;
  wire u_cosa_mux2to1_5_mux2to1_and0;
  wire u_cosa_mux2to1_5_mux2to1_not0;
  wire u_cosa_mux2to1_5_mux2to1_and1;
  wire u_cosa_mux2to1_5_mux2to1_xor0;
  wire u_cosa_mux2to1_6_mux2to1_and0;
  wire u_cosa_mux2to1_6_mux2to1_not0;
  wire u_cosa_mux2to1_6_mux2to1_and1;
  wire u_cosa_mux2to1_6_mux2to1_xor0;
  wire u_cosa_mux2to1_7_mux2to1_and0;
  wire u_cosa_mux2to1_7_mux2to1_not0;
  wire u_cosa_mux2to1_7_mux2to1_and1;
  wire u_cosa_mux2to1_7_mux2to1_xor0;
  wire u_cosa_mux2to1_8_mux2to1_and0;
  wire u_cosa_mux2to1_8_mux2to1_not0;
  wire u_cosa_mux2to1_8_mux2to1_and1;
  wire u_cosa_mux2to1_8_mux2to1_xor0;
  wire u_cosa_fa7_fa_xor0;
  wire u_cosa_fa7_fa_and0;
  wire u_cosa_fa8_fa_xor0;
  wire u_cosa_fa8_fa_and0;
  wire u_cosa_fa8_fa_xor1_not;
  wire u_cosa_fa8_fa_or0;
  wire u_cosa_mux2to1_9_mux2to1_and0;
  wire u_cosa_mux2to1_9_mux2to1_not0;
  wire u_cosa_mux2to1_9_mux2to1_and1;
  wire u_cosa_mux2to1_9_mux2to1_xor0;
  wire u_cosa_fa9_fa_xor0;
  wire u_cosa_fa9_fa_and0;
  wire u_cosa_fa10_fa_xor0;
  wire u_cosa_fa10_fa_and0;
  wire u_cosa_fa10_fa_xor1_not;
  wire u_cosa_fa10_fa_or0;
  wire u_cosa_mux2to1_10_mux2to1_and0;
  wire u_cosa_mux2to1_10_mux2to1_not0;
  wire u_cosa_mux2to1_10_mux2to1_and1;
  wire u_cosa_mux2to1_10_mux2to1_xor0;
  wire u_cosa_mux2to1_11_mux2to1_and0;
  wire u_cosa_mux2to1_11_mux2to1_not0;
  wire u_cosa_mux2to1_11_mux2to1_and1;
  wire u_cosa_mux2to1_11_mux2to1_xor0;
  wire u_cosa_mux2to1_12_mux2to1_and0;
  wire u_cosa_mux2to1_12_mux2to1_not0;
  wire u_cosa_mux2to1_12_mux2to1_and1;
  wire u_cosa_mux2to1_12_mux2to1_xor0;
  wire u_cosa_mux2to1_13_mux2to1_and0;
  wire u_cosa_mux2to1_13_mux2to1_not0;
  wire u_cosa_mux2to1_13_mux2to1_and1;
  wire u_cosa_mux2to1_13_mux2to1_xor0;
  wire u_cosa_mux2to1_14_mux2to1_and0;
  wire u_cosa_mux2to1_14_mux2to1_not0;
  wire u_cosa_mux2to1_14_mux2to1_and1;
  wire u_cosa_mux2to1_14_mux2to1_xor0;
  wire u_cosa_fa11_fa_xor0;
  wire u_cosa_fa11_fa_and0;
  wire u_cosa_fa12_fa_xor0;
  wire u_cosa_fa12_fa_and0;
  wire u_cosa_fa12_fa_xor1_not;
  wire u_cosa_fa12_fa_or0;
  wire u_cosa_mux2to1_15_mux2to1_and0;
  wire u_cosa_mux2to1_15_mux2to1_not0;
  wire u_cosa_mux2to1_15_mux2to1_and1;
  wire u_cosa_mux2to1_15_mux2to1_xor0;
  wire u_cosa_mux2to1_16_mux2to1_and0;
  wire u_cosa_mux2to1_16_mux2to1_not0;
  wire u_cosa_mux2to1_16_mux2to1_and1;
  wire u_cosa_mux2to1_16_mux2to1_xor0;
  wire u_cosa_mux2to1_17_mux2to1_and0;
  wire u_cosa_mux2to1_17_mux2to1_not0;
  wire u_cosa_mux2to1_17_mux2to1_and1;
  wire u_cosa_mux2to1_17_mux2to1_xor0;
  wire u_cosa_fa13_fa_xor0;
  wire u_cosa_fa13_fa_and0;
  wire u_cosa_fa14_fa_xor0;
  wire u_cosa_fa14_fa_and0;
  wire u_cosa_fa14_fa_xor1_not;
  wire u_cosa_fa14_fa_or0;
  wire u_cosa_mux2to1_18_mux2to1_and0;
  wire u_cosa_mux2to1_18_mux2to1_not0;
  wire u_cosa_mux2to1_18_mux2to1_and1;
  wire u_cosa_mux2to1_18_mux2to1_xor0;
  wire u_cosa_mux2to1_19_mux2to1_and0;
  wire u_cosa_mux2to1_19_mux2to1_not0;
  wire u_cosa_mux2to1_19_mux2to1_and1;
  wire u_cosa_mux2to1_19_mux2to1_xor0;
  wire u_cosa_mux2to1_20_mux2to1_and0;
  wire u_cosa_mux2to1_20_mux2to1_not0;
  wire u_cosa_mux2to1_20_mux2to1_and1;
  wire u_cosa_mux2to1_20_mux2to1_xor0;
  wire u_cosa_mux2to1_21_mux2to1_and0;
  wire u_cosa_mux2to1_21_mux2to1_not0;
  wire u_cosa_mux2to1_21_mux2to1_and1;
  wire u_cosa_mux2to1_21_mux2to1_xor0;
  wire u_cosa_mux2to1_22_mux2to1_and0;
  wire u_cosa_mux2to1_22_mux2to1_not0;
  wire u_cosa_mux2to1_22_mux2to1_and1;
  wire u_cosa_mux2to1_22_mux2to1_xor0;
  wire u_cosa_mux2to1_23_mux2to1_and0;
  wire u_cosa_mux2to1_23_mux2to1_not0;
  wire u_cosa_mux2to1_23_mux2to1_and1;
  wire u_cosa_mux2to1_23_mux2to1_xor0;
  wire u_cosa_mux2to1_24_mux2to1_and0;
  wire u_cosa_mux2to1_24_mux2to1_not0;
  wire u_cosa_mux2to1_24_mux2to1_and1;
  wire u_cosa_mux2to1_24_mux2to1_xor0;
  wire u_cosa_mux2to1_25_mux2to1_and0;
  wire u_cosa_mux2to1_25_mux2to1_not0;
  wire u_cosa_mux2to1_25_mux2to1_and1;
  wire u_cosa_mux2to1_25_mux2to1_xor0;
  wire u_cosa_mux2to1_26_mux2to1_and0;
  wire u_cosa_mux2to1_26_mux2to1_not0;
  wire u_cosa_mux2to1_26_mux2to1_and1;
  wire u_cosa_mux2to1_26_mux2to1_xor0;
  wire u_cosa_mux2to1_27_mux2to1_and0;
  wire u_cosa_mux2to1_27_mux2to1_not0;
  wire u_cosa_mux2to1_27_mux2to1_and1;
  wire u_cosa_mux2to1_27_mux2to1_xor0;

  assign u_cosa_fa0_fa_xor0 = a[0] ^ b[0];
  assign u_cosa_fa0_fa_and0 = a[0] & b[0];
  assign u_cosa_fa1_fa_xor0 = a[1] ^ b[1];
  assign u_cosa_fa1_fa_and0 = a[1] & b[1];
  assign u_cosa_fa2_fa_xor0 = a[1] ^ b[1];
  assign u_cosa_fa2_fa_and0 = a[1] & b[1];
  assign u_cosa_fa2_fa_xor1_not = ~u_cosa_fa2_fa_xor0;
  assign u_cosa_fa2_fa_or0 = u_cosa_fa2_fa_and0 | u_cosa_fa2_fa_xor0;
  assign u_cosa_mux2to1_0_mux2to1_and0 = u_cosa_fa2_fa_xor1_not & u_cosa_fa0_fa_and0;
  assign u_cosa_mux2to1_0_mux2to1_not0 = ~u_cosa_fa0_fa_and0;
  assign u_cosa_mux2to1_0_mux2to1_and1 = u_cosa_fa1_fa_xor0 & u_cosa_mux2to1_0_mux2to1_not0;
  assign u_cosa_mux2to1_0_mux2to1_xor0 = u_cosa_mux2to1_0_mux2to1_and0 ^ u_cosa_mux2to1_0_mux2to1_and1;
  assign u_cosa_mux2to1_1_mux2to1_and0 = u_cosa_fa2_fa_or0 & u_cosa_fa0_fa_and0;
  assign u_cosa_mux2to1_1_mux2to1_not0 = ~u_cosa_fa0_fa_and0;
  assign u_cosa_mux2to1_1_mux2to1_and1 = u_cosa_fa1_fa_and0 & u_cosa_mux2to1_1_mux2to1_not0;
  assign u_cosa_mux2to1_1_mux2to1_xor0 = u_cosa_mux2to1_1_mux2to1_and0 ^ u_cosa_mux2to1_1_mux2to1_and1;
  assign u_cosa_fa3_fa_xor0 = a[2] ^ b[2];
  assign u_cosa_fa3_fa_and0 = a[2] & b[2];
  assign u_cosa_fa4_fa_xor0 = a[2] ^ b[2];
  assign u_cosa_fa4_fa_and0 = a[2] & b[2];
  assign u_cosa_fa4_fa_xor1_not = ~u_cosa_fa4_fa_xor0;
  assign u_cosa_fa4_fa_or0 = u_cosa_fa4_fa_and0 | u_cosa_fa4_fa_xor0;
  assign u_cosa_mux2to1_2_mux2to1_and0 = u_cosa_fa4_fa_xor1_not & u_cosa_mux2to1_1_mux2to1_xor0;
  assign u_cosa_mux2to1_2_mux2to1_not0 = ~u_cosa_mux2to1_1_mux2to1_xor0;
  assign u_cosa_mux2to1_2_mux2to1_and1 = u_cosa_fa3_fa_xor0 & u_cosa_mux2to1_2_mux2to1_not0;
  assign u_cosa_mux2to1_2_mux2to1_xor0 = u_cosa_mux2to1_2_mux2to1_and0 ^ u_cosa_mux2to1_2_mux2to1_and1;
  assign u_cosa_fa5_fa_xor0 = a[3] ^ b[3];
  assign u_cosa_fa5_fa_and0 = a[3] & b[3];
  assign u_cosa_fa6_fa_xor0 = a[3] ^ b[3];
  assign u_cosa_fa6_fa_and0 = a[3] & b[3];
  assign u_cosa_fa6_fa_xor1_not = ~u_cosa_fa6_fa_xor0;
  assign u_cosa_fa6_fa_or0 = u_cosa_fa6_fa_and0 | u_cosa_fa6_fa_xor0;
  assign u_cosa_mux2to1_3_mux2to1_and0 = u_cosa_fa6_fa_xor1_not & u_cosa_fa3_fa_and0;
  assign u_cosa_mux2to1_3_mux2to1_not0 = ~u_cosa_fa3_fa_and0;
  assign u_cosa_mux2to1_3_mux2to1_and1 = u_cosa_fa5_fa_xor0 & u_cosa_mux2to1_3_mux2to1_not0;
  assign u_cosa_mux2to1_3_mux2to1_xor0 = u_cosa_mux2to1_3_mux2to1_and0 ^ u_cosa_mux2to1_3_mux2to1_and1;
  assign u_cosa_mux2to1_4_mux2to1_and0 = u_cosa_fa6_fa_xor1_not & u_cosa_fa4_fa_or0;
  assign u_cosa_mux2to1_4_mux2to1_not0 = ~u_cosa_fa4_fa_or0;
  assign u_cosa_mux2to1_4_mux2to1_and1 = u_cosa_fa5_fa_xor0 & u_cosa_mux2to1_4_mux2to1_not0;
  assign u_cosa_mux2to1_4_mux2to1_xor0 = u_cosa_mux2to1_4_mux2to1_and0 ^ u_cosa_mux2to1_4_mux2to1_and1;
  assign u_cosa_mux2to1_5_mux2to1_and0 = u_cosa_fa6_fa_or0 & u_cosa_fa3_fa_and0;
  assign u_cosa_mux2to1_5_mux2to1_not0 = ~u_cosa_fa3_fa_and0;
  assign u_cosa_mux2to1_5_mux2to1_and1 = u_cosa_fa5_fa_and0 & u_cosa_mux2to1_5_mux2to1_not0;
  assign u_cosa_mux2to1_5_mux2to1_xor0 = u_cosa_mux2to1_5_mux2to1_and0 ^ u_cosa_mux2to1_5_mux2to1_and1;
  assign u_cosa_mux2to1_6_mux2to1_and0 = u_cosa_fa6_fa_or0 & u_cosa_fa4_fa_or0;
  assign u_cosa_mux2to1_6_mux2to1_not0 = ~u_cosa_fa4_fa_or0;
  assign u_cosa_mux2to1_6_mux2to1_and1 = u_cosa_fa5_fa_and0 & u_cosa_mux2to1_6_mux2to1_not0;
  assign u_cosa_mux2to1_6_mux2to1_xor0 = u_cosa_mux2to1_6_mux2to1_and0 ^ u_cosa_mux2to1_6_mux2to1_and1;
  assign u_cosa_mux2to1_7_mux2to1_and0 = u_cosa_mux2to1_4_mux2to1_xor0 & u_cosa_mux2to1_1_mux2to1_xor0;
  assign u_cosa_mux2to1_7_mux2to1_not0 = ~u_cosa_mux2to1_1_mux2to1_xor0;
  assign u_cosa_mux2to1_7_mux2to1_and1 = u_cosa_mux2to1_3_mux2to1_xor0 & u_cosa_mux2to1_7_mux2to1_not0;
  assign u_cosa_mux2to1_7_mux2to1_xor0 = u_cosa_mux2to1_7_mux2to1_and0 ^ u_cosa_mux2to1_7_mux2to1_and1;
  assign u_cosa_mux2to1_8_mux2to1_and0 = u_cosa_mux2to1_6_mux2to1_xor0 & u_cosa_mux2to1_1_mux2to1_xor0;
  assign u_cosa_mux2to1_8_mux2to1_not0 = ~u_cosa_mux2to1_1_mux2to1_xor0;
  assign u_cosa_mux2to1_8_mux2to1_and1 = u_cosa_mux2to1_5_mux2to1_xor0 & u_cosa_mux2to1_8_mux2to1_not0;
  assign u_cosa_mux2to1_8_mux2to1_xor0 = u_cosa_mux2to1_8_mux2to1_and0 ^ u_cosa_mux2to1_8_mux2to1_and1;
  assign u_cosa_fa7_fa_xor0 = a[4] ^ b[4];
  assign u_cosa_fa7_fa_and0 = a[4] & b[4];
  assign u_cosa_fa8_fa_xor0 = a[4] ^ b[4];
  assign u_cosa_fa8_fa_and0 = a[4] & b[4];
  assign u_cosa_fa8_fa_xor1_not = ~u_cosa_fa8_fa_xor0;
  assign u_cosa_fa8_fa_or0 = u_cosa_fa8_fa_and0 | u_cosa_fa8_fa_xor0;
  assign u_cosa_mux2to1_9_mux2to1_and0 = u_cosa_fa8_fa_xor1_not & u_cosa_mux2to1_8_mux2to1_xor0;
  assign u_cosa_mux2to1_9_mux2to1_not0 = ~u_cosa_mux2to1_8_mux2to1_xor0;
  assign u_cosa_mux2to1_9_mux2to1_and1 = u_cosa_fa7_fa_xor0 & u_cosa_mux2to1_9_mux2to1_not0;
  assign u_cosa_mux2to1_9_mux2to1_xor0 = u_cosa_mux2to1_9_mux2to1_and0 ^ u_cosa_mux2to1_9_mux2to1_and1;
  assign u_cosa_fa9_fa_xor0 = a[5] ^ b[5];
  assign u_cosa_fa9_fa_and0 = a[5] & b[5];
  assign u_cosa_fa10_fa_xor0 = a[5] ^ b[5];
  assign u_cosa_fa10_fa_and0 = a[5] & b[5];
  assign u_cosa_fa10_fa_xor1_not = ~u_cosa_fa10_fa_xor0;
  assign u_cosa_fa10_fa_or0 = u_cosa_fa10_fa_and0 | u_cosa_fa10_fa_xor0;
  assign u_cosa_mux2to1_10_mux2to1_and0 = u_cosa_fa10_fa_xor1_not & u_cosa_fa7_fa_and0;
  assign u_cosa_mux2to1_10_mux2to1_not0 = ~u_cosa_fa7_fa_and0;
  assign u_cosa_mux2to1_10_mux2to1_and1 = u_cosa_fa9_fa_xor0 & u_cosa_mux2to1_10_mux2to1_not0;
  assign u_cosa_mux2to1_10_mux2to1_xor0 = u_cosa_mux2to1_10_mux2to1_and0 ^ u_cosa_mux2to1_10_mux2to1_and1;
  assign u_cosa_mux2to1_11_mux2to1_and0 = u_cosa_fa10_fa_xor1_not & u_cosa_fa8_fa_or0;
  assign u_cosa_mux2to1_11_mux2to1_not0 = ~u_cosa_fa8_fa_or0;
  assign u_cosa_mux2to1_11_mux2to1_and1 = u_cosa_fa9_fa_xor0 & u_cosa_mux2to1_11_mux2to1_not0;
  assign u_cosa_mux2to1_11_mux2to1_xor0 = u_cosa_mux2to1_11_mux2to1_and0 ^ u_cosa_mux2to1_11_mux2to1_and1;
  assign u_cosa_mux2to1_12_mux2to1_and0 = u_cosa_fa10_fa_or0 & u_cosa_fa7_fa_and0;
  assign u_cosa_mux2to1_12_mux2to1_not0 = ~u_cosa_fa7_fa_and0;
  assign u_cosa_mux2to1_12_mux2to1_and1 = u_cosa_fa9_fa_and0 & u_cosa_mux2to1_12_mux2to1_not0;
  assign u_cosa_mux2to1_12_mux2to1_xor0 = u_cosa_mux2to1_12_mux2to1_and0 ^ u_cosa_mux2to1_12_mux2to1_and1;
  assign u_cosa_mux2to1_13_mux2to1_and0 = u_cosa_fa10_fa_or0 & u_cosa_fa8_fa_or0;
  assign u_cosa_mux2to1_13_mux2to1_not0 = ~u_cosa_fa8_fa_or0;
  assign u_cosa_mux2to1_13_mux2to1_and1 = u_cosa_fa9_fa_and0 & u_cosa_mux2to1_13_mux2to1_not0;
  assign u_cosa_mux2to1_13_mux2to1_xor0 = u_cosa_mux2to1_13_mux2to1_and0 ^ u_cosa_mux2to1_13_mux2to1_and1;
  assign u_cosa_mux2to1_14_mux2to1_and0 = u_cosa_mux2to1_11_mux2to1_xor0 & u_cosa_mux2to1_8_mux2to1_xor0;
  assign u_cosa_mux2to1_14_mux2to1_not0 = ~u_cosa_mux2to1_8_mux2to1_xor0;
  assign u_cosa_mux2to1_14_mux2to1_and1 = u_cosa_mux2to1_10_mux2to1_xor0 & u_cosa_mux2to1_14_mux2to1_not0;
  assign u_cosa_mux2to1_14_mux2to1_xor0 = u_cosa_mux2to1_14_mux2to1_and0 ^ u_cosa_mux2to1_14_mux2to1_and1;
  assign u_cosa_fa11_fa_xor0 = a[6] ^ b[6];
  assign u_cosa_fa11_fa_and0 = a[6] & b[6];
  assign u_cosa_fa12_fa_xor0 = a[6] ^ b[6];
  assign u_cosa_fa12_fa_and0 = a[6] & b[6];
  assign u_cosa_fa12_fa_xor1_not = ~u_cosa_fa12_fa_xor0;
  assign u_cosa_fa12_fa_or0 = u_cosa_fa12_fa_and0 | u_cosa_fa12_fa_xor0;
  assign u_cosa_mux2to1_15_mux2to1_and0 = u_cosa_fa12_fa_xor1_not & u_cosa_mux2to1_12_mux2to1_xor0;
  assign u_cosa_mux2to1_15_mux2to1_not0 = ~u_cosa_mux2to1_12_mux2to1_xor0;
  assign u_cosa_mux2to1_15_mux2to1_and1 = u_cosa_fa11_fa_xor0 & u_cosa_mux2to1_15_mux2to1_not0;
  assign u_cosa_mux2to1_15_mux2to1_xor0 = u_cosa_mux2to1_15_mux2to1_and0 ^ u_cosa_mux2to1_15_mux2to1_and1;
  assign u_cosa_mux2to1_16_mux2to1_and0 = u_cosa_fa12_fa_xor1_not & u_cosa_mux2to1_13_mux2to1_xor0;
  assign u_cosa_mux2to1_16_mux2to1_not0 = ~u_cosa_mux2to1_13_mux2to1_xor0;
  assign u_cosa_mux2to1_16_mux2to1_and1 = u_cosa_mux2to1_15_mux2to1_xor0 & u_cosa_mux2to1_16_mux2to1_not0;
  assign u_cosa_mux2to1_16_mux2to1_xor0 = u_cosa_mux2to1_16_mux2to1_and0 ^ u_cosa_mux2to1_16_mux2to1_and1;
  assign u_cosa_mux2to1_17_mux2to1_and0 = u_cosa_mux2to1_16_mux2to1_xor0 & u_cosa_mux2to1_8_mux2to1_xor0;
  assign u_cosa_mux2to1_17_mux2to1_not0 = ~u_cosa_mux2to1_8_mux2to1_xor0;
  assign u_cosa_mux2to1_17_mux2to1_and1 = u_cosa_mux2to1_15_mux2to1_xor0 & u_cosa_mux2to1_17_mux2to1_not0;
  assign u_cosa_mux2to1_17_mux2to1_xor0 = u_cosa_mux2to1_17_mux2to1_and0 ^ u_cosa_mux2to1_17_mux2to1_and1;
  assign u_cosa_fa13_fa_xor0 = a[7] ^ b[7];
  assign u_cosa_fa13_fa_and0 = a[7] & b[7];
  assign u_cosa_fa14_fa_xor0 = a[7] ^ b[7];
  assign u_cosa_fa14_fa_and0 = a[7] & b[7];
  assign u_cosa_fa14_fa_xor1_not = ~u_cosa_fa14_fa_xor0;
  assign u_cosa_fa14_fa_or0 = u_cosa_fa14_fa_and0 | u_cosa_fa14_fa_xor0;
  assign u_cosa_mux2to1_18_mux2to1_and0 = u_cosa_fa14_fa_xor1_not & u_cosa_fa11_fa_and0;
  assign u_cosa_mux2to1_18_mux2to1_not0 = ~u_cosa_fa11_fa_and0;
  assign u_cosa_mux2to1_18_mux2to1_and1 = u_cosa_fa13_fa_xor0 & u_cosa_mux2to1_18_mux2to1_not0;
  assign u_cosa_mux2to1_18_mux2to1_xor0 = u_cosa_mux2to1_18_mux2to1_and0 ^ u_cosa_mux2to1_18_mux2to1_and1;
  assign u_cosa_mux2to1_19_mux2to1_and0 = u_cosa_fa14_fa_xor1_not & u_cosa_fa12_fa_or0;
  assign u_cosa_mux2to1_19_mux2to1_not0 = ~u_cosa_fa12_fa_or0;
  assign u_cosa_mux2to1_19_mux2to1_and1 = u_cosa_fa13_fa_xor0 & u_cosa_mux2to1_19_mux2to1_not0;
  assign u_cosa_mux2to1_19_mux2to1_xor0 = u_cosa_mux2to1_19_mux2to1_and0 ^ u_cosa_mux2to1_19_mux2to1_and1;
  assign u_cosa_mux2to1_20_mux2to1_and0 = u_cosa_fa14_fa_or0 & u_cosa_fa11_fa_and0;
  assign u_cosa_mux2to1_20_mux2to1_not0 = ~u_cosa_fa11_fa_and0;
  assign u_cosa_mux2to1_20_mux2to1_and1 = u_cosa_fa13_fa_and0 & u_cosa_mux2to1_20_mux2to1_not0;
  assign u_cosa_mux2to1_20_mux2to1_xor0 = u_cosa_mux2to1_20_mux2to1_and0 ^ u_cosa_mux2to1_20_mux2to1_and1;
  assign u_cosa_mux2to1_21_mux2to1_and0 = u_cosa_fa14_fa_or0 & u_cosa_fa12_fa_or0;
  assign u_cosa_mux2to1_21_mux2to1_not0 = ~u_cosa_fa12_fa_or0;
  assign u_cosa_mux2to1_21_mux2to1_and1 = u_cosa_fa13_fa_and0 & u_cosa_mux2to1_21_mux2to1_not0;
  assign u_cosa_mux2to1_21_mux2to1_xor0 = u_cosa_mux2to1_21_mux2to1_and0 ^ u_cosa_mux2to1_21_mux2to1_and1;
  assign u_cosa_mux2to1_22_mux2to1_and0 = u_cosa_mux2to1_19_mux2to1_xor0 & u_cosa_mux2to1_12_mux2to1_xor0;
  assign u_cosa_mux2to1_22_mux2to1_not0 = ~u_cosa_mux2to1_12_mux2to1_xor0;
  assign u_cosa_mux2to1_22_mux2to1_and1 = u_cosa_mux2to1_18_mux2to1_xor0 & u_cosa_mux2to1_22_mux2to1_not0;
  assign u_cosa_mux2to1_22_mux2to1_xor0 = u_cosa_mux2to1_22_mux2to1_and0 ^ u_cosa_mux2to1_22_mux2to1_and1;
  assign u_cosa_mux2to1_23_mux2to1_and0 = u_cosa_mux2to1_19_mux2to1_xor0 & u_cosa_mux2to1_13_mux2to1_xor0;
  assign u_cosa_mux2to1_23_mux2to1_not0 = ~u_cosa_mux2to1_13_mux2to1_xor0;
  assign u_cosa_mux2to1_23_mux2to1_and1 = u_cosa_mux2to1_18_mux2to1_xor0 & u_cosa_mux2to1_23_mux2to1_not0;
  assign u_cosa_mux2to1_23_mux2to1_xor0 = u_cosa_mux2to1_23_mux2to1_and0 ^ u_cosa_mux2to1_23_mux2to1_and1;
  assign u_cosa_mux2to1_24_mux2to1_and0 = u_cosa_mux2to1_21_mux2to1_xor0 & u_cosa_mux2to1_12_mux2to1_xor0;
  assign u_cosa_mux2to1_24_mux2to1_not0 = ~u_cosa_mux2to1_12_mux2to1_xor0;
  assign u_cosa_mux2to1_24_mux2to1_and1 = u_cosa_mux2to1_20_mux2to1_xor0 & u_cosa_mux2to1_24_mux2to1_not0;
  assign u_cosa_mux2to1_24_mux2to1_xor0 = u_cosa_mux2to1_24_mux2to1_and0 ^ u_cosa_mux2to1_24_mux2to1_and1;
  assign u_cosa_mux2to1_25_mux2to1_and0 = u_cosa_mux2to1_21_mux2to1_xor0 & u_cosa_mux2to1_13_mux2to1_xor0;
  assign u_cosa_mux2to1_25_mux2to1_not0 = ~u_cosa_mux2to1_13_mux2to1_xor0;
  assign u_cosa_mux2to1_25_mux2to1_and1 = u_cosa_mux2to1_20_mux2to1_xor0 & u_cosa_mux2to1_25_mux2to1_not0;
  assign u_cosa_mux2to1_25_mux2to1_xor0 = u_cosa_mux2to1_25_mux2to1_and0 ^ u_cosa_mux2to1_25_mux2to1_and1;
  assign u_cosa_mux2to1_26_mux2to1_and0 = u_cosa_mux2to1_23_mux2to1_xor0 & u_cosa_mux2to1_8_mux2to1_xor0;
  assign u_cosa_mux2to1_26_mux2to1_not0 = ~u_cosa_mux2to1_8_mux2to1_xor0;
  assign u_cosa_mux2to1_26_mux2to1_and1 = u_cosa_mux2to1_22_mux2to1_xor0 & u_cosa_mux2to1_26_mux2to1_not0;
  assign u_cosa_mux2to1_26_mux2to1_xor0 = u_cosa_mux2to1_26_mux2to1_and0 ^ u_cosa_mux2to1_26_mux2to1_and1;
  assign u_cosa_mux2to1_27_mux2to1_and0 = u_cosa_mux2to1_25_mux2to1_xor0 & u_cosa_mux2to1_8_mux2to1_xor0;
  assign u_cosa_mux2to1_27_mux2to1_not0 = ~u_cosa_mux2to1_8_mux2to1_xor0;
  assign u_cosa_mux2to1_27_mux2to1_and1 = u_cosa_mux2to1_24_mux2to1_xor0 & u_cosa_mux2to1_27_mux2to1_not0;
  assign u_cosa_mux2to1_27_mux2to1_xor0 = u_cosa_mux2to1_27_mux2to1_and0 ^ u_cosa_mux2to1_27_mux2to1_and1;

  assign u_cosa_out[0] = u_cosa_fa0_fa_xor0;
  assign u_cosa_out[1] = u_cosa_mux2to1_0_mux2to1_xor0;
  assign u_cosa_out[2] = u_cosa_mux2to1_2_mux2to1_xor0;
  assign u_cosa_out[3] = u_cosa_mux2to1_7_mux2to1_xor0;
  assign u_cosa_out[4] = u_cosa_mux2to1_9_mux2to1_xor0;
  assign u_cosa_out[5] = u_cosa_mux2to1_14_mux2to1_xor0;
  assign u_cosa_out[6] = u_cosa_mux2to1_17_mux2to1_xor0;
  assign u_cosa_out[7] = u_cosa_mux2to1_26_mux2to1_xor0;
  assign u_cosa_out[8] = u_cosa_mux2to1_27_mux2to1_xor0;
endmodule