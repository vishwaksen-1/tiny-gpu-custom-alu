module arrdiv(input [7:0] a, input [7:0] b, output [7:0] arrdiv_out);
  wire arrdiv_fs0_fs_xor0;
  wire arrdiv_fs0_fs_not0;
  wire arrdiv_fs0_fs_and0;
  wire arrdiv_fs0_fs_not1;
  wire arrdiv_fs1_fs_xor1;
  wire arrdiv_fs1_fs_not1;
  wire arrdiv_fs1_fs_and1;
  wire arrdiv_fs1_fs_or0;
  wire arrdiv_fs2_fs_xor1;
  wire arrdiv_fs2_fs_not1;
  wire arrdiv_fs2_fs_and1;
  wire arrdiv_fs2_fs_or0;
  wire arrdiv_fs3_fs_xor1;
  wire arrdiv_fs3_fs_not1;
  wire arrdiv_fs3_fs_and1;
  wire arrdiv_fs3_fs_or0;
  wire arrdiv_fs4_fs_xor1;
  wire arrdiv_fs4_fs_not1;
  wire arrdiv_fs4_fs_and1;
  wire arrdiv_fs4_fs_or0;
  wire arrdiv_fs5_fs_xor1;
  wire arrdiv_fs5_fs_not1;
  wire arrdiv_fs5_fs_and1;
  wire arrdiv_fs5_fs_or0;
  wire arrdiv_fs6_fs_xor1;
  wire arrdiv_fs6_fs_not1;
  wire arrdiv_fs6_fs_and1;
  wire arrdiv_fs6_fs_or0;
  wire arrdiv_fs7_fs_xor1;
  wire arrdiv_fs7_fs_not1;
  wire arrdiv_fs7_fs_and1;
  wire arrdiv_fs7_fs_or0;
  wire arrdiv_mux2to10_mux2to1_and0;
  wire arrdiv_mux2to10_mux2to1_not0;
  wire arrdiv_mux2to10_mux2to1_and1;
  wire arrdiv_mux2to10_mux2to1_xor0;
  wire arrdiv_mux2to11_mux2to1_not0;
  wire arrdiv_mux2to11_mux2to1_and1;
  wire arrdiv_mux2to12_mux2to1_not0;
  wire arrdiv_mux2to12_mux2to1_and1;
  wire arrdiv_mux2to13_mux2to1_not0;
  wire arrdiv_mux2to13_mux2to1_and1;
  wire arrdiv_mux2to14_mux2to1_not0;
  wire arrdiv_mux2to14_mux2to1_and1;
  wire arrdiv_mux2to15_mux2to1_not0;
  wire arrdiv_mux2to15_mux2to1_and1;
  wire arrdiv_mux2to16_mux2to1_not0;
  wire arrdiv_mux2to16_mux2to1_and1;
  wire arrdiv_not0;
  wire arrdiv_fs8_fs_xor0;
  wire arrdiv_fs8_fs_not0;
  wire arrdiv_fs8_fs_and0;
  wire arrdiv_fs8_fs_not1;
  wire arrdiv_fs9_fs_xor0;
  wire arrdiv_fs9_fs_not0;
  wire arrdiv_fs9_fs_and0;
  wire arrdiv_fs9_fs_xor1;
  wire arrdiv_fs9_fs_not1;
  wire arrdiv_fs9_fs_and1;
  wire arrdiv_fs9_fs_or0;
  wire arrdiv_fs10_fs_xor0;
  wire arrdiv_fs10_fs_not0;
  wire arrdiv_fs10_fs_and0;
  wire arrdiv_fs10_fs_xor1;
  wire arrdiv_fs10_fs_not1;
  wire arrdiv_fs10_fs_and1;
  wire arrdiv_fs10_fs_or0;
  wire arrdiv_fs11_fs_xor0;
  wire arrdiv_fs11_fs_not0;
  wire arrdiv_fs11_fs_and0;
  wire arrdiv_fs11_fs_xor1;
  wire arrdiv_fs11_fs_not1;
  wire arrdiv_fs11_fs_and1;
  wire arrdiv_fs11_fs_or0;
  wire arrdiv_fs12_fs_xor0;
  wire arrdiv_fs12_fs_not0;
  wire arrdiv_fs12_fs_and0;
  wire arrdiv_fs12_fs_xor1;
  wire arrdiv_fs12_fs_not1;
  wire arrdiv_fs12_fs_and1;
  wire arrdiv_fs12_fs_or0;
  wire arrdiv_fs13_fs_xor0;
  wire arrdiv_fs13_fs_not0;
  wire arrdiv_fs13_fs_and0;
  wire arrdiv_fs13_fs_xor1;
  wire arrdiv_fs13_fs_not1;
  wire arrdiv_fs13_fs_and1;
  wire arrdiv_fs13_fs_or0;
  wire arrdiv_fs14_fs_xor0;
  wire arrdiv_fs14_fs_not0;
  wire arrdiv_fs14_fs_and0;
  wire arrdiv_fs14_fs_xor1;
  wire arrdiv_fs14_fs_not1;
  wire arrdiv_fs14_fs_and1;
  wire arrdiv_fs14_fs_or0;
  wire arrdiv_fs15_fs_xor0;
  wire arrdiv_fs15_fs_not0;
  wire arrdiv_fs15_fs_and0;
  wire arrdiv_fs15_fs_xor1;
  wire arrdiv_fs15_fs_not1;
  wire arrdiv_fs15_fs_and1;
  wire arrdiv_fs15_fs_or0;
  wire arrdiv_mux2to17_mux2to1_and0;
  wire arrdiv_mux2to17_mux2to1_not0;
  wire arrdiv_mux2to17_mux2to1_and1;
  wire arrdiv_mux2to17_mux2to1_xor0;
  wire arrdiv_mux2to18_mux2to1_and0;
  wire arrdiv_mux2to18_mux2to1_not0;
  wire arrdiv_mux2to18_mux2to1_and1;
  wire arrdiv_mux2to18_mux2to1_xor0;
  wire arrdiv_mux2to19_mux2to1_and0;
  wire arrdiv_mux2to19_mux2to1_not0;
  wire arrdiv_mux2to19_mux2to1_and1;
  wire arrdiv_mux2to19_mux2to1_xor0;
  wire arrdiv_mux2to110_mux2to1_and0;
  wire arrdiv_mux2to110_mux2to1_not0;
  wire arrdiv_mux2to110_mux2to1_and1;
  wire arrdiv_mux2to110_mux2to1_xor0;
  wire arrdiv_mux2to111_mux2to1_and0;
  wire arrdiv_mux2to111_mux2to1_not0;
  wire arrdiv_mux2to111_mux2to1_and1;
  wire arrdiv_mux2to111_mux2to1_xor0;
  wire arrdiv_mux2to112_mux2to1_and0;
  wire arrdiv_mux2to112_mux2to1_not0;
  wire arrdiv_mux2to112_mux2to1_and1;
  wire arrdiv_mux2to112_mux2to1_xor0;
  wire arrdiv_mux2to113_mux2to1_and0;
  wire arrdiv_mux2to113_mux2to1_not0;
  wire arrdiv_mux2to113_mux2to1_and1;
  wire arrdiv_mux2to113_mux2to1_xor0;
  wire arrdiv_not1;
  wire arrdiv_fs16_fs_xor0;
  wire arrdiv_fs16_fs_not0;
  wire arrdiv_fs16_fs_and0;
  wire arrdiv_fs16_fs_not1;
  wire arrdiv_fs17_fs_xor0;
  wire arrdiv_fs17_fs_not0;
  wire arrdiv_fs17_fs_and0;
  wire arrdiv_fs17_fs_xor1;
  wire arrdiv_fs17_fs_not1;
  wire arrdiv_fs17_fs_and1;
  wire arrdiv_fs17_fs_or0;
  wire arrdiv_fs18_fs_xor0;
  wire arrdiv_fs18_fs_not0;
  wire arrdiv_fs18_fs_and0;
  wire arrdiv_fs18_fs_xor1;
  wire arrdiv_fs18_fs_not1;
  wire arrdiv_fs18_fs_and1;
  wire arrdiv_fs18_fs_or0;
  wire arrdiv_fs19_fs_xor0;
  wire arrdiv_fs19_fs_not0;
  wire arrdiv_fs19_fs_and0;
  wire arrdiv_fs19_fs_xor1;
  wire arrdiv_fs19_fs_not1;
  wire arrdiv_fs19_fs_and1;
  wire arrdiv_fs19_fs_or0;
  wire arrdiv_fs20_fs_xor0;
  wire arrdiv_fs20_fs_not0;
  wire arrdiv_fs20_fs_and0;
  wire arrdiv_fs20_fs_xor1;
  wire arrdiv_fs20_fs_not1;
  wire arrdiv_fs20_fs_and1;
  wire arrdiv_fs20_fs_or0;
  wire arrdiv_fs21_fs_xor0;
  wire arrdiv_fs21_fs_not0;
  wire arrdiv_fs21_fs_and0;
  wire arrdiv_fs21_fs_xor1;
  wire arrdiv_fs21_fs_not1;
  wire arrdiv_fs21_fs_and1;
  wire arrdiv_fs21_fs_or0;
  wire arrdiv_fs22_fs_xor0;
  wire arrdiv_fs22_fs_not0;
  wire arrdiv_fs22_fs_and0;
  wire arrdiv_fs22_fs_xor1;
  wire arrdiv_fs22_fs_not1;
  wire arrdiv_fs22_fs_and1;
  wire arrdiv_fs22_fs_or0;
  wire arrdiv_fs23_fs_xor0;
  wire arrdiv_fs23_fs_not0;
  wire arrdiv_fs23_fs_and0;
  wire arrdiv_fs23_fs_xor1;
  wire arrdiv_fs23_fs_not1;
  wire arrdiv_fs23_fs_and1;
  wire arrdiv_fs23_fs_or0;
  wire arrdiv_mux2to114_mux2to1_and0;
  wire arrdiv_mux2to114_mux2to1_not0;
  wire arrdiv_mux2to114_mux2to1_and1;
  wire arrdiv_mux2to114_mux2to1_xor0;
  wire arrdiv_mux2to115_mux2to1_and0;
  wire arrdiv_mux2to115_mux2to1_not0;
  wire arrdiv_mux2to115_mux2to1_and1;
  wire arrdiv_mux2to115_mux2to1_xor0;
  wire arrdiv_mux2to116_mux2to1_and0;
  wire arrdiv_mux2to116_mux2to1_not0;
  wire arrdiv_mux2to116_mux2to1_and1;
  wire arrdiv_mux2to116_mux2to1_xor0;
  wire arrdiv_mux2to117_mux2to1_and0;
  wire arrdiv_mux2to117_mux2to1_not0;
  wire arrdiv_mux2to117_mux2to1_and1;
  wire arrdiv_mux2to117_mux2to1_xor0;
  wire arrdiv_mux2to118_mux2to1_and0;
  wire arrdiv_mux2to118_mux2to1_not0;
  wire arrdiv_mux2to118_mux2to1_and1;
  wire arrdiv_mux2to118_mux2to1_xor0;
  wire arrdiv_mux2to119_mux2to1_and0;
  wire arrdiv_mux2to119_mux2to1_not0;
  wire arrdiv_mux2to119_mux2to1_and1;
  wire arrdiv_mux2to119_mux2to1_xor0;
  wire arrdiv_mux2to120_mux2to1_and0;
  wire arrdiv_mux2to120_mux2to1_not0;
  wire arrdiv_mux2to120_mux2to1_and1;
  wire arrdiv_mux2to120_mux2to1_xor0;
  wire arrdiv_not2;
  wire arrdiv_fs24_fs_xor0;
  wire arrdiv_fs24_fs_not0;
  wire arrdiv_fs24_fs_and0;
  wire arrdiv_fs24_fs_not1;
  wire arrdiv_fs25_fs_xor0;
  wire arrdiv_fs25_fs_not0;
  wire arrdiv_fs25_fs_and0;
  wire arrdiv_fs25_fs_xor1;
  wire arrdiv_fs25_fs_not1;
  wire arrdiv_fs25_fs_and1;
  wire arrdiv_fs25_fs_or0;
  wire arrdiv_fs26_fs_xor0;
  wire arrdiv_fs26_fs_not0;
  wire arrdiv_fs26_fs_and0;
  wire arrdiv_fs26_fs_xor1;
  wire arrdiv_fs26_fs_not1;
  wire arrdiv_fs26_fs_and1;
  wire arrdiv_fs26_fs_or0;
  wire arrdiv_fs27_fs_xor0;
  wire arrdiv_fs27_fs_not0;
  wire arrdiv_fs27_fs_and0;
  wire arrdiv_fs27_fs_xor1;
  wire arrdiv_fs27_fs_not1;
  wire arrdiv_fs27_fs_and1;
  wire arrdiv_fs27_fs_or0;
  wire arrdiv_fs28_fs_xor0;
  wire arrdiv_fs28_fs_not0;
  wire arrdiv_fs28_fs_and0;
  wire arrdiv_fs28_fs_xor1;
  wire arrdiv_fs28_fs_not1;
  wire arrdiv_fs28_fs_and1;
  wire arrdiv_fs28_fs_or0;
  wire arrdiv_fs29_fs_xor0;
  wire arrdiv_fs29_fs_not0;
  wire arrdiv_fs29_fs_and0;
  wire arrdiv_fs29_fs_xor1;
  wire arrdiv_fs29_fs_not1;
  wire arrdiv_fs29_fs_and1;
  wire arrdiv_fs29_fs_or0;
  wire arrdiv_fs30_fs_xor0;
  wire arrdiv_fs30_fs_not0;
  wire arrdiv_fs30_fs_and0;
  wire arrdiv_fs30_fs_xor1;
  wire arrdiv_fs30_fs_not1;
  wire arrdiv_fs30_fs_and1;
  wire arrdiv_fs30_fs_or0;
  wire arrdiv_fs31_fs_xor0;
  wire arrdiv_fs31_fs_not0;
  wire arrdiv_fs31_fs_and0;
  wire arrdiv_fs31_fs_xor1;
  wire arrdiv_fs31_fs_not1;
  wire arrdiv_fs31_fs_and1;
  wire arrdiv_fs31_fs_or0;
  wire arrdiv_mux2to121_mux2to1_and0;
  wire arrdiv_mux2to121_mux2to1_not0;
  wire arrdiv_mux2to121_mux2to1_and1;
  wire arrdiv_mux2to121_mux2to1_xor0;
  wire arrdiv_mux2to122_mux2to1_and0;
  wire arrdiv_mux2to122_mux2to1_not0;
  wire arrdiv_mux2to122_mux2to1_and1;
  wire arrdiv_mux2to122_mux2to1_xor0;
  wire arrdiv_mux2to123_mux2to1_and0;
  wire arrdiv_mux2to123_mux2to1_not0;
  wire arrdiv_mux2to123_mux2to1_and1;
  wire arrdiv_mux2to123_mux2to1_xor0;
  wire arrdiv_mux2to124_mux2to1_and0;
  wire arrdiv_mux2to124_mux2to1_not0;
  wire arrdiv_mux2to124_mux2to1_and1;
  wire arrdiv_mux2to124_mux2to1_xor0;
  wire arrdiv_mux2to125_mux2to1_and0;
  wire arrdiv_mux2to125_mux2to1_not0;
  wire arrdiv_mux2to125_mux2to1_and1;
  wire arrdiv_mux2to125_mux2to1_xor0;
  wire arrdiv_mux2to126_mux2to1_and0;
  wire arrdiv_mux2to126_mux2to1_not0;
  wire arrdiv_mux2to126_mux2to1_and1;
  wire arrdiv_mux2to126_mux2to1_xor0;
  wire arrdiv_mux2to127_mux2to1_and0;
  wire arrdiv_mux2to127_mux2to1_not0;
  wire arrdiv_mux2to127_mux2to1_and1;
  wire arrdiv_mux2to127_mux2to1_xor0;
  wire arrdiv_not3;
  wire arrdiv_fs32_fs_xor0;
  wire arrdiv_fs32_fs_not0;
  wire arrdiv_fs32_fs_and0;
  wire arrdiv_fs32_fs_not1;
  wire arrdiv_fs33_fs_xor0;
  wire arrdiv_fs33_fs_not0;
  wire arrdiv_fs33_fs_and0;
  wire arrdiv_fs33_fs_xor1;
  wire arrdiv_fs33_fs_not1;
  wire arrdiv_fs33_fs_and1;
  wire arrdiv_fs33_fs_or0;
  wire arrdiv_fs34_fs_xor0;
  wire arrdiv_fs34_fs_not0;
  wire arrdiv_fs34_fs_and0;
  wire arrdiv_fs34_fs_xor1;
  wire arrdiv_fs34_fs_not1;
  wire arrdiv_fs34_fs_and1;
  wire arrdiv_fs34_fs_or0;
  wire arrdiv_fs35_fs_xor0;
  wire arrdiv_fs35_fs_not0;
  wire arrdiv_fs35_fs_and0;
  wire arrdiv_fs35_fs_xor1;
  wire arrdiv_fs35_fs_not1;
  wire arrdiv_fs35_fs_and1;
  wire arrdiv_fs35_fs_or0;
  wire arrdiv_fs36_fs_xor0;
  wire arrdiv_fs36_fs_not0;
  wire arrdiv_fs36_fs_and0;
  wire arrdiv_fs36_fs_xor1;
  wire arrdiv_fs36_fs_not1;
  wire arrdiv_fs36_fs_and1;
  wire arrdiv_fs36_fs_or0;
  wire arrdiv_fs37_fs_xor0;
  wire arrdiv_fs37_fs_not0;
  wire arrdiv_fs37_fs_and0;
  wire arrdiv_fs37_fs_xor1;
  wire arrdiv_fs37_fs_not1;
  wire arrdiv_fs37_fs_and1;
  wire arrdiv_fs37_fs_or0;
  wire arrdiv_fs38_fs_xor0;
  wire arrdiv_fs38_fs_not0;
  wire arrdiv_fs38_fs_and0;
  wire arrdiv_fs38_fs_xor1;
  wire arrdiv_fs38_fs_not1;
  wire arrdiv_fs38_fs_and1;
  wire arrdiv_fs38_fs_or0;
  wire arrdiv_fs39_fs_xor0;
  wire arrdiv_fs39_fs_not0;
  wire arrdiv_fs39_fs_and0;
  wire arrdiv_fs39_fs_xor1;
  wire arrdiv_fs39_fs_not1;
  wire arrdiv_fs39_fs_and1;
  wire arrdiv_fs39_fs_or0;
  wire arrdiv_mux2to128_mux2to1_and0;
  wire arrdiv_mux2to128_mux2to1_not0;
  wire arrdiv_mux2to128_mux2to1_and1;
  wire arrdiv_mux2to128_mux2to1_xor0;
  wire arrdiv_mux2to129_mux2to1_and0;
  wire arrdiv_mux2to129_mux2to1_not0;
  wire arrdiv_mux2to129_mux2to1_and1;
  wire arrdiv_mux2to129_mux2to1_xor0;
  wire arrdiv_mux2to130_mux2to1_and0;
  wire arrdiv_mux2to130_mux2to1_not0;
  wire arrdiv_mux2to130_mux2to1_and1;
  wire arrdiv_mux2to130_mux2to1_xor0;
  wire arrdiv_mux2to131_mux2to1_and0;
  wire arrdiv_mux2to131_mux2to1_not0;
  wire arrdiv_mux2to131_mux2to1_and1;
  wire arrdiv_mux2to131_mux2to1_xor0;
  wire arrdiv_mux2to132_mux2to1_and0;
  wire arrdiv_mux2to132_mux2to1_not0;
  wire arrdiv_mux2to132_mux2to1_and1;
  wire arrdiv_mux2to132_mux2to1_xor0;
  wire arrdiv_mux2to133_mux2to1_and0;
  wire arrdiv_mux2to133_mux2to1_not0;
  wire arrdiv_mux2to133_mux2to1_and1;
  wire arrdiv_mux2to133_mux2to1_xor0;
  wire arrdiv_mux2to134_mux2to1_and0;
  wire arrdiv_mux2to134_mux2to1_not0;
  wire arrdiv_mux2to134_mux2to1_and1;
  wire arrdiv_mux2to134_mux2to1_xor0;
  wire arrdiv_not4;
  wire arrdiv_fs40_fs_xor0;
  wire arrdiv_fs40_fs_not0;
  wire arrdiv_fs40_fs_and0;
  wire arrdiv_fs40_fs_not1;
  wire arrdiv_fs41_fs_xor0;
  wire arrdiv_fs41_fs_not0;
  wire arrdiv_fs41_fs_and0;
  wire arrdiv_fs41_fs_xor1;
  wire arrdiv_fs41_fs_not1;
  wire arrdiv_fs41_fs_and1;
  wire arrdiv_fs41_fs_or0;
  wire arrdiv_fs42_fs_xor0;
  wire arrdiv_fs42_fs_not0;
  wire arrdiv_fs42_fs_and0;
  wire arrdiv_fs42_fs_xor1;
  wire arrdiv_fs42_fs_not1;
  wire arrdiv_fs42_fs_and1;
  wire arrdiv_fs42_fs_or0;
  wire arrdiv_fs43_fs_xor0;
  wire arrdiv_fs43_fs_not0;
  wire arrdiv_fs43_fs_and0;
  wire arrdiv_fs43_fs_xor1;
  wire arrdiv_fs43_fs_not1;
  wire arrdiv_fs43_fs_and1;
  wire arrdiv_fs43_fs_or0;
  wire arrdiv_fs44_fs_xor0;
  wire arrdiv_fs44_fs_not0;
  wire arrdiv_fs44_fs_and0;
  wire arrdiv_fs44_fs_xor1;
  wire arrdiv_fs44_fs_not1;
  wire arrdiv_fs44_fs_and1;
  wire arrdiv_fs44_fs_or0;
  wire arrdiv_fs45_fs_xor0;
  wire arrdiv_fs45_fs_not0;
  wire arrdiv_fs45_fs_and0;
  wire arrdiv_fs45_fs_xor1;
  wire arrdiv_fs45_fs_not1;
  wire arrdiv_fs45_fs_and1;
  wire arrdiv_fs45_fs_or0;
  wire arrdiv_fs46_fs_xor0;
  wire arrdiv_fs46_fs_not0;
  wire arrdiv_fs46_fs_and0;
  wire arrdiv_fs46_fs_xor1;
  wire arrdiv_fs46_fs_not1;
  wire arrdiv_fs46_fs_and1;
  wire arrdiv_fs46_fs_or0;
  wire arrdiv_fs47_fs_xor0;
  wire arrdiv_fs47_fs_not0;
  wire arrdiv_fs47_fs_and0;
  wire arrdiv_fs47_fs_xor1;
  wire arrdiv_fs47_fs_not1;
  wire arrdiv_fs47_fs_and1;
  wire arrdiv_fs47_fs_or0;
  wire arrdiv_mux2to135_mux2to1_and0;
  wire arrdiv_mux2to135_mux2to1_not0;
  wire arrdiv_mux2to135_mux2to1_and1;
  wire arrdiv_mux2to135_mux2to1_xor0;
  wire arrdiv_mux2to136_mux2to1_and0;
  wire arrdiv_mux2to136_mux2to1_not0;
  wire arrdiv_mux2to136_mux2to1_and1;
  wire arrdiv_mux2to136_mux2to1_xor0;
  wire arrdiv_mux2to137_mux2to1_and0;
  wire arrdiv_mux2to137_mux2to1_not0;
  wire arrdiv_mux2to137_mux2to1_and1;
  wire arrdiv_mux2to137_mux2to1_xor0;
  wire arrdiv_mux2to138_mux2to1_and0;
  wire arrdiv_mux2to138_mux2to1_not0;
  wire arrdiv_mux2to138_mux2to1_and1;
  wire arrdiv_mux2to138_mux2to1_xor0;
  wire arrdiv_mux2to139_mux2to1_and0;
  wire arrdiv_mux2to139_mux2to1_not0;
  wire arrdiv_mux2to139_mux2to1_and1;
  wire arrdiv_mux2to139_mux2to1_xor0;
  wire arrdiv_mux2to140_mux2to1_and0;
  wire arrdiv_mux2to140_mux2to1_not0;
  wire arrdiv_mux2to140_mux2to1_and1;
  wire arrdiv_mux2to140_mux2to1_xor0;
  wire arrdiv_mux2to141_mux2to1_and0;
  wire arrdiv_mux2to141_mux2to1_not0;
  wire arrdiv_mux2to141_mux2to1_and1;
  wire arrdiv_mux2to141_mux2to1_xor0;
  wire arrdiv_not5;
  wire arrdiv_fs48_fs_xor0;
  wire arrdiv_fs48_fs_not0;
  wire arrdiv_fs48_fs_and0;
  wire arrdiv_fs48_fs_not1;
  wire arrdiv_fs49_fs_xor0;
  wire arrdiv_fs49_fs_not0;
  wire arrdiv_fs49_fs_and0;
  wire arrdiv_fs49_fs_xor1;
  wire arrdiv_fs49_fs_not1;
  wire arrdiv_fs49_fs_and1;
  wire arrdiv_fs49_fs_or0;
  wire arrdiv_fs50_fs_xor0;
  wire arrdiv_fs50_fs_not0;
  wire arrdiv_fs50_fs_and0;
  wire arrdiv_fs50_fs_xor1;
  wire arrdiv_fs50_fs_not1;
  wire arrdiv_fs50_fs_and1;
  wire arrdiv_fs50_fs_or0;
  wire arrdiv_fs51_fs_xor0;
  wire arrdiv_fs51_fs_not0;
  wire arrdiv_fs51_fs_and0;
  wire arrdiv_fs51_fs_xor1;
  wire arrdiv_fs51_fs_not1;
  wire arrdiv_fs51_fs_and1;
  wire arrdiv_fs51_fs_or0;
  wire arrdiv_fs52_fs_xor0;
  wire arrdiv_fs52_fs_not0;
  wire arrdiv_fs52_fs_and0;
  wire arrdiv_fs52_fs_xor1;
  wire arrdiv_fs52_fs_not1;
  wire arrdiv_fs52_fs_and1;
  wire arrdiv_fs52_fs_or0;
  wire arrdiv_fs53_fs_xor0;
  wire arrdiv_fs53_fs_not0;
  wire arrdiv_fs53_fs_and0;
  wire arrdiv_fs53_fs_xor1;
  wire arrdiv_fs53_fs_not1;
  wire arrdiv_fs53_fs_and1;
  wire arrdiv_fs53_fs_or0;
  wire arrdiv_fs54_fs_xor0;
  wire arrdiv_fs54_fs_not0;
  wire arrdiv_fs54_fs_and0;
  wire arrdiv_fs54_fs_xor1;
  wire arrdiv_fs54_fs_not1;
  wire arrdiv_fs54_fs_and1;
  wire arrdiv_fs54_fs_or0;
  wire arrdiv_fs55_fs_xor0;
  wire arrdiv_fs55_fs_not0;
  wire arrdiv_fs55_fs_and0;
  wire arrdiv_fs55_fs_xor1;
  wire arrdiv_fs55_fs_not1;
  wire arrdiv_fs55_fs_and1;
  wire arrdiv_fs55_fs_or0;
  wire arrdiv_mux2to142_mux2to1_and0;
  wire arrdiv_mux2to142_mux2to1_not0;
  wire arrdiv_mux2to142_mux2to1_and1;
  wire arrdiv_mux2to142_mux2to1_xor0;
  wire arrdiv_mux2to143_mux2to1_and0;
  wire arrdiv_mux2to143_mux2to1_not0;
  wire arrdiv_mux2to143_mux2to1_and1;
  wire arrdiv_mux2to143_mux2to1_xor0;
  wire arrdiv_mux2to144_mux2to1_and0;
  wire arrdiv_mux2to144_mux2to1_not0;
  wire arrdiv_mux2to144_mux2to1_and1;
  wire arrdiv_mux2to144_mux2to1_xor0;
  wire arrdiv_mux2to145_mux2to1_and0;
  wire arrdiv_mux2to145_mux2to1_not0;
  wire arrdiv_mux2to145_mux2to1_and1;
  wire arrdiv_mux2to145_mux2to1_xor0;
  wire arrdiv_mux2to146_mux2to1_and0;
  wire arrdiv_mux2to146_mux2to1_not0;
  wire arrdiv_mux2to146_mux2to1_and1;
  wire arrdiv_mux2to146_mux2to1_xor0;
  wire arrdiv_mux2to147_mux2to1_and0;
  wire arrdiv_mux2to147_mux2to1_not0;
  wire arrdiv_mux2to147_mux2to1_and1;
  wire arrdiv_mux2to147_mux2to1_xor0;
  wire arrdiv_mux2to148_mux2to1_and0;
  wire arrdiv_mux2to148_mux2to1_not0;
  wire arrdiv_mux2to148_mux2to1_and1;
  wire arrdiv_mux2to148_mux2to1_xor0;
  wire arrdiv_not6;
  wire arrdiv_fs56_fs_xor0;
  wire arrdiv_fs56_fs_not0;
  wire arrdiv_fs56_fs_and0;
  wire arrdiv_fs56_fs_not1;
  wire arrdiv_fs57_fs_xor0;
  wire arrdiv_fs57_fs_not0;
  wire arrdiv_fs57_fs_and0;
  wire arrdiv_fs57_fs_xor1;
  wire arrdiv_fs57_fs_not1;
  wire arrdiv_fs57_fs_and1;
  wire arrdiv_fs57_fs_or0;
  wire arrdiv_fs58_fs_xor0;
  wire arrdiv_fs58_fs_not0;
  wire arrdiv_fs58_fs_and0;
  wire arrdiv_fs58_fs_xor1;
  wire arrdiv_fs58_fs_not1;
  wire arrdiv_fs58_fs_and1;
  wire arrdiv_fs58_fs_or0;
  wire arrdiv_fs59_fs_xor0;
  wire arrdiv_fs59_fs_not0;
  wire arrdiv_fs59_fs_and0;
  wire arrdiv_fs59_fs_xor1;
  wire arrdiv_fs59_fs_not1;
  wire arrdiv_fs59_fs_and1;
  wire arrdiv_fs59_fs_or0;
  wire arrdiv_fs60_fs_xor0;
  wire arrdiv_fs60_fs_not0;
  wire arrdiv_fs60_fs_and0;
  wire arrdiv_fs60_fs_xor1;
  wire arrdiv_fs60_fs_not1;
  wire arrdiv_fs60_fs_and1;
  wire arrdiv_fs60_fs_or0;
  wire arrdiv_fs61_fs_xor0;
  wire arrdiv_fs61_fs_not0;
  wire arrdiv_fs61_fs_and0;
  wire arrdiv_fs61_fs_xor1;
  wire arrdiv_fs61_fs_not1;
  wire arrdiv_fs61_fs_and1;
  wire arrdiv_fs61_fs_or0;
  wire arrdiv_fs62_fs_xor0;
  wire arrdiv_fs62_fs_not0;
  wire arrdiv_fs62_fs_and0;
  wire arrdiv_fs62_fs_xor1;
  wire arrdiv_fs62_fs_not1;
  wire arrdiv_fs62_fs_and1;
  wire arrdiv_fs62_fs_or0;
  wire arrdiv_fs63_fs_xor0;
  wire arrdiv_fs63_fs_not0;
  wire arrdiv_fs63_fs_and0;
  wire arrdiv_fs63_fs_xor1;
  wire arrdiv_fs63_fs_not1;
  wire arrdiv_fs63_fs_and1;
  wire arrdiv_fs63_fs_or0;
  wire arrdiv_not7;

  assign arrdiv_fs0_fs_xor0 = a[7] ^ b[0];
  assign arrdiv_fs0_fs_not0 = ~a[7];
  assign arrdiv_fs0_fs_and0 = arrdiv_fs0_fs_not0 & b[0];
  assign arrdiv_fs0_fs_not1 = ~arrdiv_fs0_fs_xor0;
  assign arrdiv_fs1_fs_xor1 = arrdiv_fs0_fs_and0 ^ b[1];
  assign arrdiv_fs1_fs_not1 = ~b[1];
  assign arrdiv_fs1_fs_and1 = arrdiv_fs1_fs_not1 & arrdiv_fs0_fs_and0;
  assign arrdiv_fs1_fs_or0 = arrdiv_fs1_fs_and1 | b[1];
  assign arrdiv_fs2_fs_xor1 = arrdiv_fs1_fs_or0 ^ b[2];
  assign arrdiv_fs2_fs_not1 = ~b[2];
  assign arrdiv_fs2_fs_and1 = arrdiv_fs2_fs_not1 & arrdiv_fs1_fs_or0;
  assign arrdiv_fs2_fs_or0 = arrdiv_fs2_fs_and1 | b[2];
  assign arrdiv_fs3_fs_xor1 = arrdiv_fs2_fs_or0 ^ b[3];
  assign arrdiv_fs3_fs_not1 = ~b[3];
  assign arrdiv_fs3_fs_and1 = arrdiv_fs3_fs_not1 & arrdiv_fs2_fs_or0;
  assign arrdiv_fs3_fs_or0 = arrdiv_fs3_fs_and1 | b[3];
  assign arrdiv_fs4_fs_xor1 = arrdiv_fs3_fs_or0 ^ b[4];
  assign arrdiv_fs4_fs_not1 = ~b[4];
  assign arrdiv_fs4_fs_and1 = arrdiv_fs4_fs_not1 & arrdiv_fs3_fs_or0;
  assign arrdiv_fs4_fs_or0 = arrdiv_fs4_fs_and1 | b[4];
  assign arrdiv_fs5_fs_xor1 = arrdiv_fs4_fs_or0 ^ b[5];
  assign arrdiv_fs5_fs_not1 = ~b[5];
  assign arrdiv_fs5_fs_and1 = arrdiv_fs5_fs_not1 & arrdiv_fs4_fs_or0;
  assign arrdiv_fs5_fs_or0 = arrdiv_fs5_fs_and1 | b[5];
  assign arrdiv_fs6_fs_xor1 = arrdiv_fs5_fs_or0 ^ b[6];
  assign arrdiv_fs6_fs_not1 = ~b[6];
  assign arrdiv_fs6_fs_and1 = arrdiv_fs6_fs_not1 & arrdiv_fs5_fs_or0;
  assign arrdiv_fs6_fs_or0 = arrdiv_fs6_fs_and1 | b[6];
  assign arrdiv_fs7_fs_xor1 = arrdiv_fs6_fs_or0 ^ b[7];
  assign arrdiv_fs7_fs_not1 = ~b[7];
  assign arrdiv_fs7_fs_and1 = arrdiv_fs7_fs_not1 & arrdiv_fs6_fs_or0;
  assign arrdiv_fs7_fs_or0 = arrdiv_fs7_fs_and1 | b[7];
  assign arrdiv_mux2to10_mux2to1_and0 = a[7] & arrdiv_fs7_fs_or0;
  assign arrdiv_mux2to10_mux2to1_not0 = ~arrdiv_fs7_fs_or0;
  assign arrdiv_mux2to10_mux2to1_and1 = arrdiv_fs0_fs_xor0 & arrdiv_mux2to10_mux2to1_not0;
  assign arrdiv_mux2to10_mux2to1_xor0 = arrdiv_mux2to10_mux2to1_and0 ^ arrdiv_mux2to10_mux2to1_and1;
  assign arrdiv_mux2to11_mux2to1_not0 = ~arrdiv_fs7_fs_or0;
  assign arrdiv_mux2to11_mux2to1_and1 = arrdiv_fs1_fs_xor1 & arrdiv_mux2to11_mux2to1_not0;
  assign arrdiv_mux2to12_mux2to1_not0 = ~arrdiv_fs7_fs_or0;
  assign arrdiv_mux2to12_mux2to1_and1 = arrdiv_fs2_fs_xor1 & arrdiv_mux2to12_mux2to1_not0;
  assign arrdiv_mux2to13_mux2to1_not0 = ~arrdiv_fs7_fs_or0;
  assign arrdiv_mux2to13_mux2to1_and1 = arrdiv_fs3_fs_xor1 & arrdiv_mux2to13_mux2to1_not0;
  assign arrdiv_mux2to14_mux2to1_not0 = ~arrdiv_fs7_fs_or0;
  assign arrdiv_mux2to14_mux2to1_and1 = arrdiv_fs4_fs_xor1 & arrdiv_mux2to14_mux2to1_not0;
  assign arrdiv_mux2to15_mux2to1_not0 = ~arrdiv_fs7_fs_or0;
  assign arrdiv_mux2to15_mux2to1_and1 = arrdiv_fs5_fs_xor1 & arrdiv_mux2to15_mux2to1_not0;
  assign arrdiv_mux2to16_mux2to1_not0 = ~arrdiv_fs7_fs_or0;
  assign arrdiv_mux2to16_mux2to1_and1 = arrdiv_fs6_fs_xor1 & arrdiv_mux2to16_mux2to1_not0;
  assign arrdiv_not0 = ~arrdiv_fs7_fs_or0;
  assign arrdiv_fs8_fs_xor0 = a[6] ^ b[0];
  assign arrdiv_fs8_fs_not0 = ~a[6];
  assign arrdiv_fs8_fs_and0 = arrdiv_fs8_fs_not0 & b[0];
  assign arrdiv_fs8_fs_not1 = ~arrdiv_fs8_fs_xor0;
  assign arrdiv_fs9_fs_xor0 = arrdiv_mux2to10_mux2to1_xor0 ^ b[1];
  assign arrdiv_fs9_fs_not0 = ~arrdiv_mux2to10_mux2to1_xor0;
  assign arrdiv_fs9_fs_and0 = arrdiv_fs9_fs_not0 & b[1];
  assign arrdiv_fs9_fs_xor1 = arrdiv_fs8_fs_and0 ^ arrdiv_fs9_fs_xor0;
  assign arrdiv_fs9_fs_not1 = ~arrdiv_fs9_fs_xor0;
  assign arrdiv_fs9_fs_and1 = arrdiv_fs9_fs_not1 & arrdiv_fs8_fs_and0;
  assign arrdiv_fs9_fs_or0 = arrdiv_fs9_fs_and1 | arrdiv_fs9_fs_and0;
  assign arrdiv_fs10_fs_xor0 = arrdiv_mux2to11_mux2to1_and1 ^ b[2];
  assign arrdiv_fs10_fs_not0 = ~arrdiv_mux2to11_mux2to1_and1;
  assign arrdiv_fs10_fs_and0 = arrdiv_fs10_fs_not0 & b[2];
  assign arrdiv_fs10_fs_xor1 = arrdiv_fs9_fs_or0 ^ arrdiv_fs10_fs_xor0;
  assign arrdiv_fs10_fs_not1 = ~arrdiv_fs10_fs_xor0;
  assign arrdiv_fs10_fs_and1 = arrdiv_fs10_fs_not1 & arrdiv_fs9_fs_or0;
  assign arrdiv_fs10_fs_or0 = arrdiv_fs10_fs_and1 | arrdiv_fs10_fs_and0;
  assign arrdiv_fs11_fs_xor0 = arrdiv_mux2to12_mux2to1_and1 ^ b[3];
  assign arrdiv_fs11_fs_not0 = ~arrdiv_mux2to12_mux2to1_and1;
  assign arrdiv_fs11_fs_and0 = arrdiv_fs11_fs_not0 & b[3];
  assign arrdiv_fs11_fs_xor1 = arrdiv_fs10_fs_or0 ^ arrdiv_fs11_fs_xor0;
  assign arrdiv_fs11_fs_not1 = ~arrdiv_fs11_fs_xor0;
  assign arrdiv_fs11_fs_and1 = arrdiv_fs11_fs_not1 & arrdiv_fs10_fs_or0;
  assign arrdiv_fs11_fs_or0 = arrdiv_fs11_fs_and1 | arrdiv_fs11_fs_and0;
  assign arrdiv_fs12_fs_xor0 = arrdiv_mux2to13_mux2to1_and1 ^ b[4];
  assign arrdiv_fs12_fs_not0 = ~arrdiv_mux2to13_mux2to1_and1;
  assign arrdiv_fs12_fs_and0 = arrdiv_fs12_fs_not0 & b[4];
  assign arrdiv_fs12_fs_xor1 = arrdiv_fs11_fs_or0 ^ arrdiv_fs12_fs_xor0;
  assign arrdiv_fs12_fs_not1 = ~arrdiv_fs12_fs_xor0;
  assign arrdiv_fs12_fs_and1 = arrdiv_fs12_fs_not1 & arrdiv_fs11_fs_or0;
  assign arrdiv_fs12_fs_or0 = arrdiv_fs12_fs_and1 | arrdiv_fs12_fs_and0;
  assign arrdiv_fs13_fs_xor0 = arrdiv_mux2to14_mux2to1_and1 ^ b[5];
  assign arrdiv_fs13_fs_not0 = ~arrdiv_mux2to14_mux2to1_and1;
  assign arrdiv_fs13_fs_and0 = arrdiv_fs13_fs_not0 & b[5];
  assign arrdiv_fs13_fs_xor1 = arrdiv_fs12_fs_or0 ^ arrdiv_fs13_fs_xor0;
  assign arrdiv_fs13_fs_not1 = ~arrdiv_fs13_fs_xor0;
  assign arrdiv_fs13_fs_and1 = arrdiv_fs13_fs_not1 & arrdiv_fs12_fs_or0;
  assign arrdiv_fs13_fs_or0 = arrdiv_fs13_fs_and1 | arrdiv_fs13_fs_and0;
  assign arrdiv_fs14_fs_xor0 = arrdiv_mux2to15_mux2to1_and1 ^ b[6];
  assign arrdiv_fs14_fs_not0 = ~arrdiv_mux2to15_mux2to1_and1;
  assign arrdiv_fs14_fs_and0 = arrdiv_fs14_fs_not0 & b[6];
  assign arrdiv_fs14_fs_xor1 = arrdiv_fs13_fs_or0 ^ arrdiv_fs14_fs_xor0;
  assign arrdiv_fs14_fs_not1 = ~arrdiv_fs14_fs_xor0;
  assign arrdiv_fs14_fs_and1 = arrdiv_fs14_fs_not1 & arrdiv_fs13_fs_or0;
  assign arrdiv_fs14_fs_or0 = arrdiv_fs14_fs_and1 | arrdiv_fs14_fs_and0;
  assign arrdiv_fs15_fs_xor0 = arrdiv_mux2to16_mux2to1_and1 ^ b[7];
  assign arrdiv_fs15_fs_not0 = ~arrdiv_mux2to16_mux2to1_and1;
  assign arrdiv_fs15_fs_and0 = arrdiv_fs15_fs_not0 & b[7];
  assign arrdiv_fs15_fs_xor1 = arrdiv_fs14_fs_or0 ^ arrdiv_fs15_fs_xor0;
  assign arrdiv_fs15_fs_not1 = ~arrdiv_fs15_fs_xor0;
  assign arrdiv_fs15_fs_and1 = arrdiv_fs15_fs_not1 & arrdiv_fs14_fs_or0;
  assign arrdiv_fs15_fs_or0 = arrdiv_fs15_fs_and1 | arrdiv_fs15_fs_and0;
  assign arrdiv_mux2to17_mux2to1_and0 = a[6] & arrdiv_fs15_fs_or0;
  assign arrdiv_mux2to17_mux2to1_not0 = ~arrdiv_fs15_fs_or0;
  assign arrdiv_mux2to17_mux2to1_and1 = arrdiv_fs8_fs_xor0 & arrdiv_mux2to17_mux2to1_not0;
  assign arrdiv_mux2to17_mux2to1_xor0 = arrdiv_mux2to17_mux2to1_and0 ^ arrdiv_mux2to17_mux2to1_and1;
  assign arrdiv_mux2to18_mux2to1_and0 = arrdiv_mux2to10_mux2to1_xor0 & arrdiv_fs15_fs_or0;
  assign arrdiv_mux2to18_mux2to1_not0 = ~arrdiv_fs15_fs_or0;
  assign arrdiv_mux2to18_mux2to1_and1 = arrdiv_fs9_fs_xor1 & arrdiv_mux2to18_mux2to1_not0;
  assign arrdiv_mux2to18_mux2to1_xor0 = arrdiv_mux2to18_mux2to1_and0 ^ arrdiv_mux2to18_mux2to1_and1;
  assign arrdiv_mux2to19_mux2to1_and0 = arrdiv_mux2to11_mux2to1_and1 & arrdiv_fs15_fs_or0;
  assign arrdiv_mux2to19_mux2to1_not0 = ~arrdiv_fs15_fs_or0;
  assign arrdiv_mux2to19_mux2to1_and1 = arrdiv_fs10_fs_xor1 & arrdiv_mux2to19_mux2to1_not0;
  assign arrdiv_mux2to19_mux2to1_xor0 = arrdiv_mux2to19_mux2to1_and0 ^ arrdiv_mux2to19_mux2to1_and1;
  assign arrdiv_mux2to110_mux2to1_and0 = arrdiv_mux2to12_mux2to1_and1 & arrdiv_fs15_fs_or0;
  assign arrdiv_mux2to110_mux2to1_not0 = ~arrdiv_fs15_fs_or0;
  assign arrdiv_mux2to110_mux2to1_and1 = arrdiv_fs11_fs_xor1 & arrdiv_mux2to110_mux2to1_not0;
  assign arrdiv_mux2to110_mux2to1_xor0 = arrdiv_mux2to110_mux2to1_and0 ^ arrdiv_mux2to110_mux2to1_and1;
  assign arrdiv_mux2to111_mux2to1_and0 = arrdiv_mux2to13_mux2to1_and1 & arrdiv_fs15_fs_or0;
  assign arrdiv_mux2to111_mux2to1_not0 = ~arrdiv_fs15_fs_or0;
  assign arrdiv_mux2to111_mux2to1_and1 = arrdiv_fs12_fs_xor1 & arrdiv_mux2to111_mux2to1_not0;
  assign arrdiv_mux2to111_mux2to1_xor0 = arrdiv_mux2to111_mux2to1_and0 ^ arrdiv_mux2to111_mux2to1_and1;
  assign arrdiv_mux2to112_mux2to1_and0 = arrdiv_mux2to14_mux2to1_and1 & arrdiv_fs15_fs_or0;
  assign arrdiv_mux2to112_mux2to1_not0 = ~arrdiv_fs15_fs_or0;
  assign arrdiv_mux2to112_mux2to1_and1 = arrdiv_fs13_fs_xor1 & arrdiv_mux2to112_mux2to1_not0;
  assign arrdiv_mux2to112_mux2to1_xor0 = arrdiv_mux2to112_mux2to1_and0 ^ arrdiv_mux2to112_mux2to1_and1;
  assign arrdiv_mux2to113_mux2to1_and0 = arrdiv_mux2to15_mux2to1_and1 & arrdiv_fs15_fs_or0;
  assign arrdiv_mux2to113_mux2to1_not0 = ~arrdiv_fs15_fs_or0;
  assign arrdiv_mux2to113_mux2to1_and1 = arrdiv_fs14_fs_xor1 & arrdiv_mux2to113_mux2to1_not0;
  assign arrdiv_mux2to113_mux2to1_xor0 = arrdiv_mux2to113_mux2to1_and0 ^ arrdiv_mux2to113_mux2to1_and1;
  assign arrdiv_not1 = ~arrdiv_fs15_fs_or0;
  assign arrdiv_fs16_fs_xor0 = a[5] ^ b[0];
  assign arrdiv_fs16_fs_not0 = ~a[5];
  assign arrdiv_fs16_fs_and0 = arrdiv_fs16_fs_not0 & b[0];
  assign arrdiv_fs16_fs_not1 = ~arrdiv_fs16_fs_xor0;
  assign arrdiv_fs17_fs_xor0 = arrdiv_mux2to17_mux2to1_xor0 ^ b[1];
  assign arrdiv_fs17_fs_not0 = ~arrdiv_mux2to17_mux2to1_xor0;
  assign arrdiv_fs17_fs_and0 = arrdiv_fs17_fs_not0 & b[1];
  assign arrdiv_fs17_fs_xor1 = arrdiv_fs16_fs_and0 ^ arrdiv_fs17_fs_xor0;
  assign arrdiv_fs17_fs_not1 = ~arrdiv_fs17_fs_xor0;
  assign arrdiv_fs17_fs_and1 = arrdiv_fs17_fs_not1 & arrdiv_fs16_fs_and0;
  assign arrdiv_fs17_fs_or0 = arrdiv_fs17_fs_and1 | arrdiv_fs17_fs_and0;
  assign arrdiv_fs18_fs_xor0 = arrdiv_mux2to18_mux2to1_xor0 ^ b[2];
  assign arrdiv_fs18_fs_not0 = ~arrdiv_mux2to18_mux2to1_xor0;
  assign arrdiv_fs18_fs_and0 = arrdiv_fs18_fs_not0 & b[2];
  assign arrdiv_fs18_fs_xor1 = arrdiv_fs17_fs_or0 ^ arrdiv_fs18_fs_xor0;
  assign arrdiv_fs18_fs_not1 = ~arrdiv_fs18_fs_xor0;
  assign arrdiv_fs18_fs_and1 = arrdiv_fs18_fs_not1 & arrdiv_fs17_fs_or0;
  assign arrdiv_fs18_fs_or0 = arrdiv_fs18_fs_and1 | arrdiv_fs18_fs_and0;
  assign arrdiv_fs19_fs_xor0 = arrdiv_mux2to19_mux2to1_xor0 ^ b[3];
  assign arrdiv_fs19_fs_not0 = ~arrdiv_mux2to19_mux2to1_xor0;
  assign arrdiv_fs19_fs_and0 = arrdiv_fs19_fs_not0 & b[3];
  assign arrdiv_fs19_fs_xor1 = arrdiv_fs18_fs_or0 ^ arrdiv_fs19_fs_xor0;
  assign arrdiv_fs19_fs_not1 = ~arrdiv_fs19_fs_xor0;
  assign arrdiv_fs19_fs_and1 = arrdiv_fs19_fs_not1 & arrdiv_fs18_fs_or0;
  assign arrdiv_fs19_fs_or0 = arrdiv_fs19_fs_and1 | arrdiv_fs19_fs_and0;
  assign arrdiv_fs20_fs_xor0 = arrdiv_mux2to110_mux2to1_xor0 ^ b[4];
  assign arrdiv_fs20_fs_not0 = ~arrdiv_mux2to110_mux2to1_xor0;
  assign arrdiv_fs20_fs_and0 = arrdiv_fs20_fs_not0 & b[4];
  assign arrdiv_fs20_fs_xor1 = arrdiv_fs19_fs_or0 ^ arrdiv_fs20_fs_xor0;
  assign arrdiv_fs20_fs_not1 = ~arrdiv_fs20_fs_xor0;
  assign arrdiv_fs20_fs_and1 = arrdiv_fs20_fs_not1 & arrdiv_fs19_fs_or0;
  assign arrdiv_fs20_fs_or0 = arrdiv_fs20_fs_and1 | arrdiv_fs20_fs_and0;
  assign arrdiv_fs21_fs_xor0 = arrdiv_mux2to111_mux2to1_xor0 ^ b[5];
  assign arrdiv_fs21_fs_not0 = ~arrdiv_mux2to111_mux2to1_xor0;
  assign arrdiv_fs21_fs_and0 = arrdiv_fs21_fs_not0 & b[5];
  assign arrdiv_fs21_fs_xor1 = arrdiv_fs20_fs_or0 ^ arrdiv_fs21_fs_xor0;
  assign arrdiv_fs21_fs_not1 = ~arrdiv_fs21_fs_xor0;
  assign arrdiv_fs21_fs_and1 = arrdiv_fs21_fs_not1 & arrdiv_fs20_fs_or0;
  assign arrdiv_fs21_fs_or0 = arrdiv_fs21_fs_and1 | arrdiv_fs21_fs_and0;
  assign arrdiv_fs22_fs_xor0 = arrdiv_mux2to112_mux2to1_xor0 ^ b[6];
  assign arrdiv_fs22_fs_not0 = ~arrdiv_mux2to112_mux2to1_xor0;
  assign arrdiv_fs22_fs_and0 = arrdiv_fs22_fs_not0 & b[6];
  assign arrdiv_fs22_fs_xor1 = arrdiv_fs21_fs_or0 ^ arrdiv_fs22_fs_xor0;
  assign arrdiv_fs22_fs_not1 = ~arrdiv_fs22_fs_xor0;
  assign arrdiv_fs22_fs_and1 = arrdiv_fs22_fs_not1 & arrdiv_fs21_fs_or0;
  assign arrdiv_fs22_fs_or0 = arrdiv_fs22_fs_and1 | arrdiv_fs22_fs_and0;
  assign arrdiv_fs23_fs_xor0 = arrdiv_mux2to113_mux2to1_xor0 ^ b[7];
  assign arrdiv_fs23_fs_not0 = ~arrdiv_mux2to113_mux2to1_xor0;
  assign arrdiv_fs23_fs_and0 = arrdiv_fs23_fs_not0 & b[7];
  assign arrdiv_fs23_fs_xor1 = arrdiv_fs22_fs_or0 ^ arrdiv_fs23_fs_xor0;
  assign arrdiv_fs23_fs_not1 = ~arrdiv_fs23_fs_xor0;
  assign arrdiv_fs23_fs_and1 = arrdiv_fs23_fs_not1 & arrdiv_fs22_fs_or0;
  assign arrdiv_fs23_fs_or0 = arrdiv_fs23_fs_and1 | arrdiv_fs23_fs_and0;
  assign arrdiv_mux2to114_mux2to1_and0 = a[5] & arrdiv_fs23_fs_or0;
  assign arrdiv_mux2to114_mux2to1_not0 = ~arrdiv_fs23_fs_or0;
  assign arrdiv_mux2to114_mux2to1_and1 = arrdiv_fs16_fs_xor0 & arrdiv_mux2to114_mux2to1_not0;
  assign arrdiv_mux2to114_mux2to1_xor0 = arrdiv_mux2to114_mux2to1_and0 ^ arrdiv_mux2to114_mux2to1_and1;
  assign arrdiv_mux2to115_mux2to1_and0 = arrdiv_mux2to17_mux2to1_xor0 & arrdiv_fs23_fs_or0;
  assign arrdiv_mux2to115_mux2to1_not0 = ~arrdiv_fs23_fs_or0;
  assign arrdiv_mux2to115_mux2to1_and1 = arrdiv_fs17_fs_xor1 & arrdiv_mux2to115_mux2to1_not0;
  assign arrdiv_mux2to115_mux2to1_xor0 = arrdiv_mux2to115_mux2to1_and0 ^ arrdiv_mux2to115_mux2to1_and1;
  assign arrdiv_mux2to116_mux2to1_and0 = arrdiv_mux2to18_mux2to1_xor0 & arrdiv_fs23_fs_or0;
  assign arrdiv_mux2to116_mux2to1_not0 = ~arrdiv_fs23_fs_or0;
  assign arrdiv_mux2to116_mux2to1_and1 = arrdiv_fs18_fs_xor1 & arrdiv_mux2to116_mux2to1_not0;
  assign arrdiv_mux2to116_mux2to1_xor0 = arrdiv_mux2to116_mux2to1_and0 ^ arrdiv_mux2to116_mux2to1_and1;
  assign arrdiv_mux2to117_mux2to1_and0 = arrdiv_mux2to19_mux2to1_xor0 & arrdiv_fs23_fs_or0;
  assign arrdiv_mux2to117_mux2to1_not0 = ~arrdiv_fs23_fs_or0;
  assign arrdiv_mux2to117_mux2to1_and1 = arrdiv_fs19_fs_xor1 & arrdiv_mux2to117_mux2to1_not0;
  assign arrdiv_mux2to117_mux2to1_xor0 = arrdiv_mux2to117_mux2to1_and0 ^ arrdiv_mux2to117_mux2to1_and1;
  assign arrdiv_mux2to118_mux2to1_and0 = arrdiv_mux2to110_mux2to1_xor0 & arrdiv_fs23_fs_or0;
  assign arrdiv_mux2to118_mux2to1_not0 = ~arrdiv_fs23_fs_or0;
  assign arrdiv_mux2to118_mux2to1_and1 = arrdiv_fs20_fs_xor1 & arrdiv_mux2to118_mux2to1_not0;
  assign arrdiv_mux2to118_mux2to1_xor0 = arrdiv_mux2to118_mux2to1_and0 ^ arrdiv_mux2to118_mux2to1_and1;
  assign arrdiv_mux2to119_mux2to1_and0 = arrdiv_mux2to111_mux2to1_xor0 & arrdiv_fs23_fs_or0;
  assign arrdiv_mux2to119_mux2to1_not0 = ~arrdiv_fs23_fs_or0;
  assign arrdiv_mux2to119_mux2to1_and1 = arrdiv_fs21_fs_xor1 & arrdiv_mux2to119_mux2to1_not0;
  assign arrdiv_mux2to119_mux2to1_xor0 = arrdiv_mux2to119_mux2to1_and0 ^ arrdiv_mux2to119_mux2to1_and1;
  assign arrdiv_mux2to120_mux2to1_and0 = arrdiv_mux2to112_mux2to1_xor0 & arrdiv_fs23_fs_or0;
  assign arrdiv_mux2to120_mux2to1_not0 = ~arrdiv_fs23_fs_or0;
  assign arrdiv_mux2to120_mux2to1_and1 = arrdiv_fs22_fs_xor1 & arrdiv_mux2to120_mux2to1_not0;
  assign arrdiv_mux2to120_mux2to1_xor0 = arrdiv_mux2to120_mux2to1_and0 ^ arrdiv_mux2to120_mux2to1_and1;
  assign arrdiv_not2 = ~arrdiv_fs23_fs_or0;
  assign arrdiv_fs24_fs_xor0 = a[4] ^ b[0];
  assign arrdiv_fs24_fs_not0 = ~a[4];
  assign arrdiv_fs24_fs_and0 = arrdiv_fs24_fs_not0 & b[0];
  assign arrdiv_fs24_fs_not1 = ~arrdiv_fs24_fs_xor0;
  assign arrdiv_fs25_fs_xor0 = arrdiv_mux2to114_mux2to1_xor0 ^ b[1];
  assign arrdiv_fs25_fs_not0 = ~arrdiv_mux2to114_mux2to1_xor0;
  assign arrdiv_fs25_fs_and0 = arrdiv_fs25_fs_not0 & b[1];
  assign arrdiv_fs25_fs_xor1 = arrdiv_fs24_fs_and0 ^ arrdiv_fs25_fs_xor0;
  assign arrdiv_fs25_fs_not1 = ~arrdiv_fs25_fs_xor0;
  assign arrdiv_fs25_fs_and1 = arrdiv_fs25_fs_not1 & arrdiv_fs24_fs_and0;
  assign arrdiv_fs25_fs_or0 = arrdiv_fs25_fs_and1 | arrdiv_fs25_fs_and0;
  assign arrdiv_fs26_fs_xor0 = arrdiv_mux2to115_mux2to1_xor0 ^ b[2];
  assign arrdiv_fs26_fs_not0 = ~arrdiv_mux2to115_mux2to1_xor0;
  assign arrdiv_fs26_fs_and0 = arrdiv_fs26_fs_not0 & b[2];
  assign arrdiv_fs26_fs_xor1 = arrdiv_fs25_fs_or0 ^ arrdiv_fs26_fs_xor0;
  assign arrdiv_fs26_fs_not1 = ~arrdiv_fs26_fs_xor0;
  assign arrdiv_fs26_fs_and1 = arrdiv_fs26_fs_not1 & arrdiv_fs25_fs_or0;
  assign arrdiv_fs26_fs_or0 = arrdiv_fs26_fs_and1 | arrdiv_fs26_fs_and0;
  assign arrdiv_fs27_fs_xor0 = arrdiv_mux2to116_mux2to1_xor0 ^ b[3];
  assign arrdiv_fs27_fs_not0 = ~arrdiv_mux2to116_mux2to1_xor0;
  assign arrdiv_fs27_fs_and0 = arrdiv_fs27_fs_not0 & b[3];
  assign arrdiv_fs27_fs_xor1 = arrdiv_fs26_fs_or0 ^ arrdiv_fs27_fs_xor0;
  assign arrdiv_fs27_fs_not1 = ~arrdiv_fs27_fs_xor0;
  assign arrdiv_fs27_fs_and1 = arrdiv_fs27_fs_not1 & arrdiv_fs26_fs_or0;
  assign arrdiv_fs27_fs_or0 = arrdiv_fs27_fs_and1 | arrdiv_fs27_fs_and0;
  assign arrdiv_fs28_fs_xor0 = arrdiv_mux2to117_mux2to1_xor0 ^ b[4];
  assign arrdiv_fs28_fs_not0 = ~arrdiv_mux2to117_mux2to1_xor0;
  assign arrdiv_fs28_fs_and0 = arrdiv_fs28_fs_not0 & b[4];
  assign arrdiv_fs28_fs_xor1 = arrdiv_fs27_fs_or0 ^ arrdiv_fs28_fs_xor0;
  assign arrdiv_fs28_fs_not1 = ~arrdiv_fs28_fs_xor0;
  assign arrdiv_fs28_fs_and1 = arrdiv_fs28_fs_not1 & arrdiv_fs27_fs_or0;
  assign arrdiv_fs28_fs_or0 = arrdiv_fs28_fs_and1 | arrdiv_fs28_fs_and0;
  assign arrdiv_fs29_fs_xor0 = arrdiv_mux2to118_mux2to1_xor0 ^ b[5];
  assign arrdiv_fs29_fs_not0 = ~arrdiv_mux2to118_mux2to1_xor0;
  assign arrdiv_fs29_fs_and0 = arrdiv_fs29_fs_not0 & b[5];
  assign arrdiv_fs29_fs_xor1 = arrdiv_fs28_fs_or0 ^ arrdiv_fs29_fs_xor0;
  assign arrdiv_fs29_fs_not1 = ~arrdiv_fs29_fs_xor0;
  assign arrdiv_fs29_fs_and1 = arrdiv_fs29_fs_not1 & arrdiv_fs28_fs_or0;
  assign arrdiv_fs29_fs_or0 = arrdiv_fs29_fs_and1 | arrdiv_fs29_fs_and0;
  assign arrdiv_fs30_fs_xor0 = arrdiv_mux2to119_mux2to1_xor0 ^ b[6];
  assign arrdiv_fs30_fs_not0 = ~arrdiv_mux2to119_mux2to1_xor0;
  assign arrdiv_fs30_fs_and0 = arrdiv_fs30_fs_not0 & b[6];
  assign arrdiv_fs30_fs_xor1 = arrdiv_fs29_fs_or0 ^ arrdiv_fs30_fs_xor0;
  assign arrdiv_fs30_fs_not1 = ~arrdiv_fs30_fs_xor0;
  assign arrdiv_fs30_fs_and1 = arrdiv_fs30_fs_not1 & arrdiv_fs29_fs_or0;
  assign arrdiv_fs30_fs_or0 = arrdiv_fs30_fs_and1 | arrdiv_fs30_fs_and0;
  assign arrdiv_fs31_fs_xor0 = arrdiv_mux2to120_mux2to1_xor0 ^ b[7];
  assign arrdiv_fs31_fs_not0 = ~arrdiv_mux2to120_mux2to1_xor0;
  assign arrdiv_fs31_fs_and0 = arrdiv_fs31_fs_not0 & b[7];
  assign arrdiv_fs31_fs_xor1 = arrdiv_fs30_fs_or0 ^ arrdiv_fs31_fs_xor0;
  assign arrdiv_fs31_fs_not1 = ~arrdiv_fs31_fs_xor0;
  assign arrdiv_fs31_fs_and1 = arrdiv_fs31_fs_not1 & arrdiv_fs30_fs_or0;
  assign arrdiv_fs31_fs_or0 = arrdiv_fs31_fs_and1 | arrdiv_fs31_fs_and0;
  assign arrdiv_mux2to121_mux2to1_and0 = a[4] & arrdiv_fs31_fs_or0;
  assign arrdiv_mux2to121_mux2to1_not0 = ~arrdiv_fs31_fs_or0;
  assign arrdiv_mux2to121_mux2to1_and1 = arrdiv_fs24_fs_xor0 & arrdiv_mux2to121_mux2to1_not0;
  assign arrdiv_mux2to121_mux2to1_xor0 = arrdiv_mux2to121_mux2to1_and0 ^ arrdiv_mux2to121_mux2to1_and1;
  assign arrdiv_mux2to122_mux2to1_and0 = arrdiv_mux2to114_mux2to1_xor0 & arrdiv_fs31_fs_or0;
  assign arrdiv_mux2to122_mux2to1_not0 = ~arrdiv_fs31_fs_or0;
  assign arrdiv_mux2to122_mux2to1_and1 = arrdiv_fs25_fs_xor1 & arrdiv_mux2to122_mux2to1_not0;
  assign arrdiv_mux2to122_mux2to1_xor0 = arrdiv_mux2to122_mux2to1_and0 ^ arrdiv_mux2to122_mux2to1_and1;
  assign arrdiv_mux2to123_mux2to1_and0 = arrdiv_mux2to115_mux2to1_xor0 & arrdiv_fs31_fs_or0;
  assign arrdiv_mux2to123_mux2to1_not0 = ~arrdiv_fs31_fs_or0;
  assign arrdiv_mux2to123_mux2to1_and1 = arrdiv_fs26_fs_xor1 & arrdiv_mux2to123_mux2to1_not0;
  assign arrdiv_mux2to123_mux2to1_xor0 = arrdiv_mux2to123_mux2to1_and0 ^ arrdiv_mux2to123_mux2to1_and1;
  assign arrdiv_mux2to124_mux2to1_and0 = arrdiv_mux2to116_mux2to1_xor0 & arrdiv_fs31_fs_or0;
  assign arrdiv_mux2to124_mux2to1_not0 = ~arrdiv_fs31_fs_or0;
  assign arrdiv_mux2to124_mux2to1_and1 = arrdiv_fs27_fs_xor1 & arrdiv_mux2to124_mux2to1_not0;
  assign arrdiv_mux2to124_mux2to1_xor0 = arrdiv_mux2to124_mux2to1_and0 ^ arrdiv_mux2to124_mux2to1_and1;
  assign arrdiv_mux2to125_mux2to1_and0 = arrdiv_mux2to117_mux2to1_xor0 & arrdiv_fs31_fs_or0;
  assign arrdiv_mux2to125_mux2to1_not0 = ~arrdiv_fs31_fs_or0;
  assign arrdiv_mux2to125_mux2to1_and1 = arrdiv_fs28_fs_xor1 & arrdiv_mux2to125_mux2to1_not0;
  assign arrdiv_mux2to125_mux2to1_xor0 = arrdiv_mux2to125_mux2to1_and0 ^ arrdiv_mux2to125_mux2to1_and1;
  assign arrdiv_mux2to126_mux2to1_and0 = arrdiv_mux2to118_mux2to1_xor0 & arrdiv_fs31_fs_or0;
  assign arrdiv_mux2to126_mux2to1_not0 = ~arrdiv_fs31_fs_or0;
  assign arrdiv_mux2to126_mux2to1_and1 = arrdiv_fs29_fs_xor1 & arrdiv_mux2to126_mux2to1_not0;
  assign arrdiv_mux2to126_mux2to1_xor0 = arrdiv_mux2to126_mux2to1_and0 ^ arrdiv_mux2to126_mux2to1_and1;
  assign arrdiv_mux2to127_mux2to1_and0 = arrdiv_mux2to119_mux2to1_xor0 & arrdiv_fs31_fs_or0;
  assign arrdiv_mux2to127_mux2to1_not0 = ~arrdiv_fs31_fs_or0;
  assign arrdiv_mux2to127_mux2to1_and1 = arrdiv_fs30_fs_xor1 & arrdiv_mux2to127_mux2to1_not0;
  assign arrdiv_mux2to127_mux2to1_xor0 = arrdiv_mux2to127_mux2to1_and0 ^ arrdiv_mux2to127_mux2to1_and1;
  assign arrdiv_not3 = ~arrdiv_fs31_fs_or0;
  assign arrdiv_fs32_fs_xor0 = a[3] ^ b[0];
  assign arrdiv_fs32_fs_not0 = ~a[3];
  assign arrdiv_fs32_fs_and0 = arrdiv_fs32_fs_not0 & b[0];
  assign arrdiv_fs32_fs_not1 = ~arrdiv_fs32_fs_xor0;
  assign arrdiv_fs33_fs_xor0 = arrdiv_mux2to121_mux2to1_xor0 ^ b[1];
  assign arrdiv_fs33_fs_not0 = ~arrdiv_mux2to121_mux2to1_xor0;
  assign arrdiv_fs33_fs_and0 = arrdiv_fs33_fs_not0 & b[1];
  assign arrdiv_fs33_fs_xor1 = arrdiv_fs32_fs_and0 ^ arrdiv_fs33_fs_xor0;
  assign arrdiv_fs33_fs_not1 = ~arrdiv_fs33_fs_xor0;
  assign arrdiv_fs33_fs_and1 = arrdiv_fs33_fs_not1 & arrdiv_fs32_fs_and0;
  assign arrdiv_fs33_fs_or0 = arrdiv_fs33_fs_and1 | arrdiv_fs33_fs_and0;
  assign arrdiv_fs34_fs_xor0 = arrdiv_mux2to122_mux2to1_xor0 ^ b[2];
  assign arrdiv_fs34_fs_not0 = ~arrdiv_mux2to122_mux2to1_xor0;
  assign arrdiv_fs34_fs_and0 = arrdiv_fs34_fs_not0 & b[2];
  assign arrdiv_fs34_fs_xor1 = arrdiv_fs33_fs_or0 ^ arrdiv_fs34_fs_xor0;
  assign arrdiv_fs34_fs_not1 = ~arrdiv_fs34_fs_xor0;
  assign arrdiv_fs34_fs_and1 = arrdiv_fs34_fs_not1 & arrdiv_fs33_fs_or0;
  assign arrdiv_fs34_fs_or0 = arrdiv_fs34_fs_and1 | arrdiv_fs34_fs_and0;
  assign arrdiv_fs35_fs_xor0 = arrdiv_mux2to123_mux2to1_xor0 ^ b[3];
  assign arrdiv_fs35_fs_not0 = ~arrdiv_mux2to123_mux2to1_xor0;
  assign arrdiv_fs35_fs_and0 = arrdiv_fs35_fs_not0 & b[3];
  assign arrdiv_fs35_fs_xor1 = arrdiv_fs34_fs_or0 ^ arrdiv_fs35_fs_xor0;
  assign arrdiv_fs35_fs_not1 = ~arrdiv_fs35_fs_xor0;
  assign arrdiv_fs35_fs_and1 = arrdiv_fs35_fs_not1 & arrdiv_fs34_fs_or0;
  assign arrdiv_fs35_fs_or0 = arrdiv_fs35_fs_and1 | arrdiv_fs35_fs_and0;
  assign arrdiv_fs36_fs_xor0 = arrdiv_mux2to124_mux2to1_xor0 ^ b[4];
  assign arrdiv_fs36_fs_not0 = ~arrdiv_mux2to124_mux2to1_xor0;
  assign arrdiv_fs36_fs_and0 = arrdiv_fs36_fs_not0 & b[4];
  assign arrdiv_fs36_fs_xor1 = arrdiv_fs35_fs_or0 ^ arrdiv_fs36_fs_xor0;
  assign arrdiv_fs36_fs_not1 = ~arrdiv_fs36_fs_xor0;
  assign arrdiv_fs36_fs_and1 = arrdiv_fs36_fs_not1 & arrdiv_fs35_fs_or0;
  assign arrdiv_fs36_fs_or0 = arrdiv_fs36_fs_and1 | arrdiv_fs36_fs_and0;
  assign arrdiv_fs37_fs_xor0 = arrdiv_mux2to125_mux2to1_xor0 ^ b[5];
  assign arrdiv_fs37_fs_not0 = ~arrdiv_mux2to125_mux2to1_xor0;
  assign arrdiv_fs37_fs_and0 = arrdiv_fs37_fs_not0 & b[5];
  assign arrdiv_fs37_fs_xor1 = arrdiv_fs36_fs_or0 ^ arrdiv_fs37_fs_xor0;
  assign arrdiv_fs37_fs_not1 = ~arrdiv_fs37_fs_xor0;
  assign arrdiv_fs37_fs_and1 = arrdiv_fs37_fs_not1 & arrdiv_fs36_fs_or0;
  assign arrdiv_fs37_fs_or0 = arrdiv_fs37_fs_and1 | arrdiv_fs37_fs_and0;
  assign arrdiv_fs38_fs_xor0 = arrdiv_mux2to126_mux2to1_xor0 ^ b[6];
  assign arrdiv_fs38_fs_not0 = ~arrdiv_mux2to126_mux2to1_xor0;
  assign arrdiv_fs38_fs_and0 = arrdiv_fs38_fs_not0 & b[6];
  assign arrdiv_fs38_fs_xor1 = arrdiv_fs37_fs_or0 ^ arrdiv_fs38_fs_xor0;
  assign arrdiv_fs38_fs_not1 = ~arrdiv_fs38_fs_xor0;
  assign arrdiv_fs38_fs_and1 = arrdiv_fs38_fs_not1 & arrdiv_fs37_fs_or0;
  assign arrdiv_fs38_fs_or0 = arrdiv_fs38_fs_and1 | arrdiv_fs38_fs_and0;
  assign arrdiv_fs39_fs_xor0 = arrdiv_mux2to127_mux2to1_xor0 ^ b[7];
  assign arrdiv_fs39_fs_not0 = ~arrdiv_mux2to127_mux2to1_xor0;
  assign arrdiv_fs39_fs_and0 = arrdiv_fs39_fs_not0 & b[7];
  assign arrdiv_fs39_fs_xor1 = arrdiv_fs38_fs_or0 ^ arrdiv_fs39_fs_xor0;
  assign arrdiv_fs39_fs_not1 = ~arrdiv_fs39_fs_xor0;
  assign arrdiv_fs39_fs_and1 = arrdiv_fs39_fs_not1 & arrdiv_fs38_fs_or0;
  assign arrdiv_fs39_fs_or0 = arrdiv_fs39_fs_and1 | arrdiv_fs39_fs_and0;
  assign arrdiv_mux2to128_mux2to1_and0 = a[3] & arrdiv_fs39_fs_or0;
  assign arrdiv_mux2to128_mux2to1_not0 = ~arrdiv_fs39_fs_or0;
  assign arrdiv_mux2to128_mux2to1_and1 = arrdiv_fs32_fs_xor0 & arrdiv_mux2to128_mux2to1_not0;
  assign arrdiv_mux2to128_mux2to1_xor0 = arrdiv_mux2to128_mux2to1_and0 ^ arrdiv_mux2to128_mux2to1_and1;
  assign arrdiv_mux2to129_mux2to1_and0 = arrdiv_mux2to121_mux2to1_xor0 & arrdiv_fs39_fs_or0;
  assign arrdiv_mux2to129_mux2to1_not0 = ~arrdiv_fs39_fs_or0;
  assign arrdiv_mux2to129_mux2to1_and1 = arrdiv_fs33_fs_xor1 & arrdiv_mux2to129_mux2to1_not0;
  assign arrdiv_mux2to129_mux2to1_xor0 = arrdiv_mux2to129_mux2to1_and0 ^ arrdiv_mux2to129_mux2to1_and1;
  assign arrdiv_mux2to130_mux2to1_and0 = arrdiv_mux2to122_mux2to1_xor0 & arrdiv_fs39_fs_or0;
  assign arrdiv_mux2to130_mux2to1_not0 = ~arrdiv_fs39_fs_or0;
  assign arrdiv_mux2to130_mux2to1_and1 = arrdiv_fs34_fs_xor1 & arrdiv_mux2to130_mux2to1_not0;
  assign arrdiv_mux2to130_mux2to1_xor0 = arrdiv_mux2to130_mux2to1_and0 ^ arrdiv_mux2to130_mux2to1_and1;
  assign arrdiv_mux2to131_mux2to1_and0 = arrdiv_mux2to123_mux2to1_xor0 & arrdiv_fs39_fs_or0;
  assign arrdiv_mux2to131_mux2to1_not0 = ~arrdiv_fs39_fs_or0;
  assign arrdiv_mux2to131_mux2to1_and1 = arrdiv_fs35_fs_xor1 & arrdiv_mux2to131_mux2to1_not0;
  assign arrdiv_mux2to131_mux2to1_xor0 = arrdiv_mux2to131_mux2to1_and0 ^ arrdiv_mux2to131_mux2to1_and1;
  assign arrdiv_mux2to132_mux2to1_and0 = arrdiv_mux2to124_mux2to1_xor0 & arrdiv_fs39_fs_or0;
  assign arrdiv_mux2to132_mux2to1_not0 = ~arrdiv_fs39_fs_or0;
  assign arrdiv_mux2to132_mux2to1_and1 = arrdiv_fs36_fs_xor1 & arrdiv_mux2to132_mux2to1_not0;
  assign arrdiv_mux2to132_mux2to1_xor0 = arrdiv_mux2to132_mux2to1_and0 ^ arrdiv_mux2to132_mux2to1_and1;
  assign arrdiv_mux2to133_mux2to1_and0 = arrdiv_mux2to125_mux2to1_xor0 & arrdiv_fs39_fs_or0;
  assign arrdiv_mux2to133_mux2to1_not0 = ~arrdiv_fs39_fs_or0;
  assign arrdiv_mux2to133_mux2to1_and1 = arrdiv_fs37_fs_xor1 & arrdiv_mux2to133_mux2to1_not0;
  assign arrdiv_mux2to133_mux2to1_xor0 = arrdiv_mux2to133_mux2to1_and0 ^ arrdiv_mux2to133_mux2to1_and1;
  assign arrdiv_mux2to134_mux2to1_and0 = arrdiv_mux2to126_mux2to1_xor0 & arrdiv_fs39_fs_or0;
  assign arrdiv_mux2to134_mux2to1_not0 = ~arrdiv_fs39_fs_or0;
  assign arrdiv_mux2to134_mux2to1_and1 = arrdiv_fs38_fs_xor1 & arrdiv_mux2to134_mux2to1_not0;
  assign arrdiv_mux2to134_mux2to1_xor0 = arrdiv_mux2to134_mux2to1_and0 ^ arrdiv_mux2to134_mux2to1_and1;
  assign arrdiv_not4 = ~arrdiv_fs39_fs_or0;
  assign arrdiv_fs40_fs_xor0 = a[2] ^ b[0];
  assign arrdiv_fs40_fs_not0 = ~a[2];
  assign arrdiv_fs40_fs_and0 = arrdiv_fs40_fs_not0 & b[0];
  assign arrdiv_fs40_fs_not1 = ~arrdiv_fs40_fs_xor0;
  assign arrdiv_fs41_fs_xor0 = arrdiv_mux2to128_mux2to1_xor0 ^ b[1];
  assign arrdiv_fs41_fs_not0 = ~arrdiv_mux2to128_mux2to1_xor0;
  assign arrdiv_fs41_fs_and0 = arrdiv_fs41_fs_not0 & b[1];
  assign arrdiv_fs41_fs_xor1 = arrdiv_fs40_fs_and0 ^ arrdiv_fs41_fs_xor0;
  assign arrdiv_fs41_fs_not1 = ~arrdiv_fs41_fs_xor0;
  assign arrdiv_fs41_fs_and1 = arrdiv_fs41_fs_not1 & arrdiv_fs40_fs_and0;
  assign arrdiv_fs41_fs_or0 = arrdiv_fs41_fs_and1 | arrdiv_fs41_fs_and0;
  assign arrdiv_fs42_fs_xor0 = arrdiv_mux2to129_mux2to1_xor0 ^ b[2];
  assign arrdiv_fs42_fs_not0 = ~arrdiv_mux2to129_mux2to1_xor0;
  assign arrdiv_fs42_fs_and0 = arrdiv_fs42_fs_not0 & b[2];
  assign arrdiv_fs42_fs_xor1 = arrdiv_fs41_fs_or0 ^ arrdiv_fs42_fs_xor0;
  assign arrdiv_fs42_fs_not1 = ~arrdiv_fs42_fs_xor0;
  assign arrdiv_fs42_fs_and1 = arrdiv_fs42_fs_not1 & arrdiv_fs41_fs_or0;
  assign arrdiv_fs42_fs_or0 = arrdiv_fs42_fs_and1 | arrdiv_fs42_fs_and0;
  assign arrdiv_fs43_fs_xor0 = arrdiv_mux2to130_mux2to1_xor0 ^ b[3];
  assign arrdiv_fs43_fs_not0 = ~arrdiv_mux2to130_mux2to1_xor0;
  assign arrdiv_fs43_fs_and0 = arrdiv_fs43_fs_not0 & b[3];
  assign arrdiv_fs43_fs_xor1 = arrdiv_fs42_fs_or0 ^ arrdiv_fs43_fs_xor0;
  assign arrdiv_fs43_fs_not1 = ~arrdiv_fs43_fs_xor0;
  assign arrdiv_fs43_fs_and1 = arrdiv_fs43_fs_not1 & arrdiv_fs42_fs_or0;
  assign arrdiv_fs43_fs_or0 = arrdiv_fs43_fs_and1 | arrdiv_fs43_fs_and0;
  assign arrdiv_fs44_fs_xor0 = arrdiv_mux2to131_mux2to1_xor0 ^ b[4];
  assign arrdiv_fs44_fs_not0 = ~arrdiv_mux2to131_mux2to1_xor0;
  assign arrdiv_fs44_fs_and0 = arrdiv_fs44_fs_not0 & b[4];
  assign arrdiv_fs44_fs_xor1 = arrdiv_fs43_fs_or0 ^ arrdiv_fs44_fs_xor0;
  assign arrdiv_fs44_fs_not1 = ~arrdiv_fs44_fs_xor0;
  assign arrdiv_fs44_fs_and1 = arrdiv_fs44_fs_not1 & arrdiv_fs43_fs_or0;
  assign arrdiv_fs44_fs_or0 = arrdiv_fs44_fs_and1 | arrdiv_fs44_fs_and0;
  assign arrdiv_fs45_fs_xor0 = arrdiv_mux2to132_mux2to1_xor0 ^ b[5];
  assign arrdiv_fs45_fs_not0 = ~arrdiv_mux2to132_mux2to1_xor0;
  assign arrdiv_fs45_fs_and0 = arrdiv_fs45_fs_not0 & b[5];
  assign arrdiv_fs45_fs_xor1 = arrdiv_fs44_fs_or0 ^ arrdiv_fs45_fs_xor0;
  assign arrdiv_fs45_fs_not1 = ~arrdiv_fs45_fs_xor0;
  assign arrdiv_fs45_fs_and1 = arrdiv_fs45_fs_not1 & arrdiv_fs44_fs_or0;
  assign arrdiv_fs45_fs_or0 = arrdiv_fs45_fs_and1 | arrdiv_fs45_fs_and0;
  assign arrdiv_fs46_fs_xor0 = arrdiv_mux2to133_mux2to1_xor0 ^ b[6];
  assign arrdiv_fs46_fs_not0 = ~arrdiv_mux2to133_mux2to1_xor0;
  assign arrdiv_fs46_fs_and0 = arrdiv_fs46_fs_not0 & b[6];
  assign arrdiv_fs46_fs_xor1 = arrdiv_fs45_fs_or0 ^ arrdiv_fs46_fs_xor0;
  assign arrdiv_fs46_fs_not1 = ~arrdiv_fs46_fs_xor0;
  assign arrdiv_fs46_fs_and1 = arrdiv_fs46_fs_not1 & arrdiv_fs45_fs_or0;
  assign arrdiv_fs46_fs_or0 = arrdiv_fs46_fs_and1 | arrdiv_fs46_fs_and0;
  assign arrdiv_fs47_fs_xor0 = arrdiv_mux2to134_mux2to1_xor0 ^ b[7];
  assign arrdiv_fs47_fs_not0 = ~arrdiv_mux2to134_mux2to1_xor0;
  assign arrdiv_fs47_fs_and0 = arrdiv_fs47_fs_not0 & b[7];
  assign arrdiv_fs47_fs_xor1 = arrdiv_fs46_fs_or0 ^ arrdiv_fs47_fs_xor0;
  assign arrdiv_fs47_fs_not1 = ~arrdiv_fs47_fs_xor0;
  assign arrdiv_fs47_fs_and1 = arrdiv_fs47_fs_not1 & arrdiv_fs46_fs_or0;
  assign arrdiv_fs47_fs_or0 = arrdiv_fs47_fs_and1 | arrdiv_fs47_fs_and0;
  assign arrdiv_mux2to135_mux2to1_and0 = a[2] & arrdiv_fs47_fs_or0;
  assign arrdiv_mux2to135_mux2to1_not0 = ~arrdiv_fs47_fs_or0;
  assign arrdiv_mux2to135_mux2to1_and1 = arrdiv_fs40_fs_xor0 & arrdiv_mux2to135_mux2to1_not0;
  assign arrdiv_mux2to135_mux2to1_xor0 = arrdiv_mux2to135_mux2to1_and0 ^ arrdiv_mux2to135_mux2to1_and1;
  assign arrdiv_mux2to136_mux2to1_and0 = arrdiv_mux2to128_mux2to1_xor0 & arrdiv_fs47_fs_or0;
  assign arrdiv_mux2to136_mux2to1_not0 = ~arrdiv_fs47_fs_or0;
  assign arrdiv_mux2to136_mux2to1_and1 = arrdiv_fs41_fs_xor1 & arrdiv_mux2to136_mux2to1_not0;
  assign arrdiv_mux2to136_mux2to1_xor0 = arrdiv_mux2to136_mux2to1_and0 ^ arrdiv_mux2to136_mux2to1_and1;
  assign arrdiv_mux2to137_mux2to1_and0 = arrdiv_mux2to129_mux2to1_xor0 & arrdiv_fs47_fs_or0;
  assign arrdiv_mux2to137_mux2to1_not0 = ~arrdiv_fs47_fs_or0;
  assign arrdiv_mux2to137_mux2to1_and1 = arrdiv_fs42_fs_xor1 & arrdiv_mux2to137_mux2to1_not0;
  assign arrdiv_mux2to137_mux2to1_xor0 = arrdiv_mux2to137_mux2to1_and0 ^ arrdiv_mux2to137_mux2to1_and1;
  assign arrdiv_mux2to138_mux2to1_and0 = arrdiv_mux2to130_mux2to1_xor0 & arrdiv_fs47_fs_or0;
  assign arrdiv_mux2to138_mux2to1_not0 = ~arrdiv_fs47_fs_or0;
  assign arrdiv_mux2to138_mux2to1_and1 = arrdiv_fs43_fs_xor1 & arrdiv_mux2to138_mux2to1_not0;
  assign arrdiv_mux2to138_mux2to1_xor0 = arrdiv_mux2to138_mux2to1_and0 ^ arrdiv_mux2to138_mux2to1_and1;
  assign arrdiv_mux2to139_mux2to1_and0 = arrdiv_mux2to131_mux2to1_xor0 & arrdiv_fs47_fs_or0;
  assign arrdiv_mux2to139_mux2to1_not0 = ~arrdiv_fs47_fs_or0;
  assign arrdiv_mux2to139_mux2to1_and1 = arrdiv_fs44_fs_xor1 & arrdiv_mux2to139_mux2to1_not0;
  assign arrdiv_mux2to139_mux2to1_xor0 = arrdiv_mux2to139_mux2to1_and0 ^ arrdiv_mux2to139_mux2to1_and1;
  assign arrdiv_mux2to140_mux2to1_and0 = arrdiv_mux2to132_mux2to1_xor0 & arrdiv_fs47_fs_or0;
  assign arrdiv_mux2to140_mux2to1_not0 = ~arrdiv_fs47_fs_or0;
  assign arrdiv_mux2to140_mux2to1_and1 = arrdiv_fs45_fs_xor1 & arrdiv_mux2to140_mux2to1_not0;
  assign arrdiv_mux2to140_mux2to1_xor0 = arrdiv_mux2to140_mux2to1_and0 ^ arrdiv_mux2to140_mux2to1_and1;
  assign arrdiv_mux2to141_mux2to1_and0 = arrdiv_mux2to133_mux2to1_xor0 & arrdiv_fs47_fs_or0;
  assign arrdiv_mux2to141_mux2to1_not0 = ~arrdiv_fs47_fs_or0;
  assign arrdiv_mux2to141_mux2to1_and1 = arrdiv_fs46_fs_xor1 & arrdiv_mux2to141_mux2to1_not0;
  assign arrdiv_mux2to141_mux2to1_xor0 = arrdiv_mux2to141_mux2to1_and0 ^ arrdiv_mux2to141_mux2to1_and1;
  assign arrdiv_not5 = ~arrdiv_fs47_fs_or0;
  assign arrdiv_fs48_fs_xor0 = a[1] ^ b[0];
  assign arrdiv_fs48_fs_not0 = ~a[1];
  assign arrdiv_fs48_fs_and0 = arrdiv_fs48_fs_not0 & b[0];
  assign arrdiv_fs48_fs_not1 = ~arrdiv_fs48_fs_xor0;
  assign arrdiv_fs49_fs_xor0 = arrdiv_mux2to135_mux2to1_xor0 ^ b[1];
  assign arrdiv_fs49_fs_not0 = ~arrdiv_mux2to135_mux2to1_xor0;
  assign arrdiv_fs49_fs_and0 = arrdiv_fs49_fs_not0 & b[1];
  assign arrdiv_fs49_fs_xor1 = arrdiv_fs48_fs_and0 ^ arrdiv_fs49_fs_xor0;
  assign arrdiv_fs49_fs_not1 = ~arrdiv_fs49_fs_xor0;
  assign arrdiv_fs49_fs_and1 = arrdiv_fs49_fs_not1 & arrdiv_fs48_fs_and0;
  assign arrdiv_fs49_fs_or0 = arrdiv_fs49_fs_and1 | arrdiv_fs49_fs_and0;
  assign arrdiv_fs50_fs_xor0 = arrdiv_mux2to136_mux2to1_xor0 ^ b[2];
  assign arrdiv_fs50_fs_not0 = ~arrdiv_mux2to136_mux2to1_xor0;
  assign arrdiv_fs50_fs_and0 = arrdiv_fs50_fs_not0 & b[2];
  assign arrdiv_fs50_fs_xor1 = arrdiv_fs49_fs_or0 ^ arrdiv_fs50_fs_xor0;
  assign arrdiv_fs50_fs_not1 = ~arrdiv_fs50_fs_xor0;
  assign arrdiv_fs50_fs_and1 = arrdiv_fs50_fs_not1 & arrdiv_fs49_fs_or0;
  assign arrdiv_fs50_fs_or0 = arrdiv_fs50_fs_and1 | arrdiv_fs50_fs_and0;
  assign arrdiv_fs51_fs_xor0 = arrdiv_mux2to137_mux2to1_xor0 ^ b[3];
  assign arrdiv_fs51_fs_not0 = ~arrdiv_mux2to137_mux2to1_xor0;
  assign arrdiv_fs51_fs_and0 = arrdiv_fs51_fs_not0 & b[3];
  assign arrdiv_fs51_fs_xor1 = arrdiv_fs50_fs_or0 ^ arrdiv_fs51_fs_xor0;
  assign arrdiv_fs51_fs_not1 = ~arrdiv_fs51_fs_xor0;
  assign arrdiv_fs51_fs_and1 = arrdiv_fs51_fs_not1 & arrdiv_fs50_fs_or0;
  assign arrdiv_fs51_fs_or0 = arrdiv_fs51_fs_and1 | arrdiv_fs51_fs_and0;
  assign arrdiv_fs52_fs_xor0 = arrdiv_mux2to138_mux2to1_xor0 ^ b[4];
  assign arrdiv_fs52_fs_not0 = ~arrdiv_mux2to138_mux2to1_xor0;
  assign arrdiv_fs52_fs_and0 = arrdiv_fs52_fs_not0 & b[4];
  assign arrdiv_fs52_fs_xor1 = arrdiv_fs51_fs_or0 ^ arrdiv_fs52_fs_xor0;
  assign arrdiv_fs52_fs_not1 = ~arrdiv_fs52_fs_xor0;
  assign arrdiv_fs52_fs_and1 = arrdiv_fs52_fs_not1 & arrdiv_fs51_fs_or0;
  assign arrdiv_fs52_fs_or0 = arrdiv_fs52_fs_and1 | arrdiv_fs52_fs_and0;
  assign arrdiv_fs53_fs_xor0 = arrdiv_mux2to139_mux2to1_xor0 ^ b[5];
  assign arrdiv_fs53_fs_not0 = ~arrdiv_mux2to139_mux2to1_xor0;
  assign arrdiv_fs53_fs_and0 = arrdiv_fs53_fs_not0 & b[5];
  assign arrdiv_fs53_fs_xor1 = arrdiv_fs52_fs_or0 ^ arrdiv_fs53_fs_xor0;
  assign arrdiv_fs53_fs_not1 = ~arrdiv_fs53_fs_xor0;
  assign arrdiv_fs53_fs_and1 = arrdiv_fs53_fs_not1 & arrdiv_fs52_fs_or0;
  assign arrdiv_fs53_fs_or0 = arrdiv_fs53_fs_and1 | arrdiv_fs53_fs_and0;
  assign arrdiv_fs54_fs_xor0 = arrdiv_mux2to140_mux2to1_xor0 ^ b[6];
  assign arrdiv_fs54_fs_not0 = ~arrdiv_mux2to140_mux2to1_xor0;
  assign arrdiv_fs54_fs_and0 = arrdiv_fs54_fs_not0 & b[6];
  assign arrdiv_fs54_fs_xor1 = arrdiv_fs53_fs_or0 ^ arrdiv_fs54_fs_xor0;
  assign arrdiv_fs54_fs_not1 = ~arrdiv_fs54_fs_xor0;
  assign arrdiv_fs54_fs_and1 = arrdiv_fs54_fs_not1 & arrdiv_fs53_fs_or0;
  assign arrdiv_fs54_fs_or0 = arrdiv_fs54_fs_and1 | arrdiv_fs54_fs_and0;
  assign arrdiv_fs55_fs_xor0 = arrdiv_mux2to141_mux2to1_xor0 ^ b[7];
  assign arrdiv_fs55_fs_not0 = ~arrdiv_mux2to141_mux2to1_xor0;
  assign arrdiv_fs55_fs_and0 = arrdiv_fs55_fs_not0 & b[7];
  assign arrdiv_fs55_fs_xor1 = arrdiv_fs54_fs_or0 ^ arrdiv_fs55_fs_xor0;
  assign arrdiv_fs55_fs_not1 = ~arrdiv_fs55_fs_xor0;
  assign arrdiv_fs55_fs_and1 = arrdiv_fs55_fs_not1 & arrdiv_fs54_fs_or0;
  assign arrdiv_fs55_fs_or0 = arrdiv_fs55_fs_and1 | arrdiv_fs55_fs_and0;
  assign arrdiv_mux2to142_mux2to1_and0 = a[1] & arrdiv_fs55_fs_or0;
  assign arrdiv_mux2to142_mux2to1_not0 = ~arrdiv_fs55_fs_or0;
  assign arrdiv_mux2to142_mux2to1_and1 = arrdiv_fs48_fs_xor0 & arrdiv_mux2to142_mux2to1_not0;
  assign arrdiv_mux2to142_mux2to1_xor0 = arrdiv_mux2to142_mux2to1_and0 ^ arrdiv_mux2to142_mux2to1_and1;
  assign arrdiv_mux2to143_mux2to1_and0 = arrdiv_mux2to135_mux2to1_xor0 & arrdiv_fs55_fs_or0;
  assign arrdiv_mux2to143_mux2to1_not0 = ~arrdiv_fs55_fs_or0;
  assign arrdiv_mux2to143_mux2to1_and1 = arrdiv_fs49_fs_xor1 & arrdiv_mux2to143_mux2to1_not0;
  assign arrdiv_mux2to143_mux2to1_xor0 = arrdiv_mux2to143_mux2to1_and0 ^ arrdiv_mux2to143_mux2to1_and1;
  assign arrdiv_mux2to144_mux2to1_and0 = arrdiv_mux2to136_mux2to1_xor0 & arrdiv_fs55_fs_or0;
  assign arrdiv_mux2to144_mux2to1_not0 = ~arrdiv_fs55_fs_or0;
  assign arrdiv_mux2to144_mux2to1_and1 = arrdiv_fs50_fs_xor1 & arrdiv_mux2to144_mux2to1_not0;
  assign arrdiv_mux2to144_mux2to1_xor0 = arrdiv_mux2to144_mux2to1_and0 ^ arrdiv_mux2to144_mux2to1_and1;
  assign arrdiv_mux2to145_mux2to1_and0 = arrdiv_mux2to137_mux2to1_xor0 & arrdiv_fs55_fs_or0;
  assign arrdiv_mux2to145_mux2to1_not0 = ~arrdiv_fs55_fs_or0;
  assign arrdiv_mux2to145_mux2to1_and1 = arrdiv_fs51_fs_xor1 & arrdiv_mux2to145_mux2to1_not0;
  assign arrdiv_mux2to145_mux2to1_xor0 = arrdiv_mux2to145_mux2to1_and0 ^ arrdiv_mux2to145_mux2to1_and1;
  assign arrdiv_mux2to146_mux2to1_and0 = arrdiv_mux2to138_mux2to1_xor0 & arrdiv_fs55_fs_or0;
  assign arrdiv_mux2to146_mux2to1_not0 = ~arrdiv_fs55_fs_or0;
  assign arrdiv_mux2to146_mux2to1_and1 = arrdiv_fs52_fs_xor1 & arrdiv_mux2to146_mux2to1_not0;
  assign arrdiv_mux2to146_mux2to1_xor0 = arrdiv_mux2to146_mux2to1_and0 ^ arrdiv_mux2to146_mux2to1_and1;
  assign arrdiv_mux2to147_mux2to1_and0 = arrdiv_mux2to139_mux2to1_xor0 & arrdiv_fs55_fs_or0;
  assign arrdiv_mux2to147_mux2to1_not0 = ~arrdiv_fs55_fs_or0;
  assign arrdiv_mux2to147_mux2to1_and1 = arrdiv_fs53_fs_xor1 & arrdiv_mux2to147_mux2to1_not0;
  assign arrdiv_mux2to147_mux2to1_xor0 = arrdiv_mux2to147_mux2to1_and0 ^ arrdiv_mux2to147_mux2to1_and1;
  assign arrdiv_mux2to148_mux2to1_and0 = arrdiv_mux2to140_mux2to1_xor0 & arrdiv_fs55_fs_or0;
  assign arrdiv_mux2to148_mux2to1_not0 = ~arrdiv_fs55_fs_or0;
  assign arrdiv_mux2to148_mux2to1_and1 = arrdiv_fs54_fs_xor1 & arrdiv_mux2to148_mux2to1_not0;
  assign arrdiv_mux2to148_mux2to1_xor0 = arrdiv_mux2to148_mux2to1_and0 ^ arrdiv_mux2to148_mux2to1_and1;
  assign arrdiv_not6 = ~arrdiv_fs55_fs_or0;
  assign arrdiv_fs56_fs_xor0 = a[0] ^ b[0];
  assign arrdiv_fs56_fs_not0 = ~a[0];
  assign arrdiv_fs56_fs_and0 = arrdiv_fs56_fs_not0 & b[0];
  assign arrdiv_fs56_fs_not1 = ~arrdiv_fs56_fs_xor0;
  assign arrdiv_fs57_fs_xor0 = arrdiv_mux2to142_mux2to1_xor0 ^ b[1];
  assign arrdiv_fs57_fs_not0 = ~arrdiv_mux2to142_mux2to1_xor0;
  assign arrdiv_fs57_fs_and0 = arrdiv_fs57_fs_not0 & b[1];
  assign arrdiv_fs57_fs_xor1 = arrdiv_fs56_fs_and0 ^ arrdiv_fs57_fs_xor0;
  assign arrdiv_fs57_fs_not1 = ~arrdiv_fs57_fs_xor0;
  assign arrdiv_fs57_fs_and1 = arrdiv_fs57_fs_not1 & arrdiv_fs56_fs_and0;
  assign arrdiv_fs57_fs_or0 = arrdiv_fs57_fs_and1 | arrdiv_fs57_fs_and0;
  assign arrdiv_fs58_fs_xor0 = arrdiv_mux2to143_mux2to1_xor0 ^ b[2];
  assign arrdiv_fs58_fs_not0 = ~arrdiv_mux2to143_mux2to1_xor0;
  assign arrdiv_fs58_fs_and0 = arrdiv_fs58_fs_not0 & b[2];
  assign arrdiv_fs58_fs_xor1 = arrdiv_fs57_fs_or0 ^ arrdiv_fs58_fs_xor0;
  assign arrdiv_fs58_fs_not1 = ~arrdiv_fs58_fs_xor0;
  assign arrdiv_fs58_fs_and1 = arrdiv_fs58_fs_not1 & arrdiv_fs57_fs_or0;
  assign arrdiv_fs58_fs_or0 = arrdiv_fs58_fs_and1 | arrdiv_fs58_fs_and0;
  assign arrdiv_fs59_fs_xor0 = arrdiv_mux2to144_mux2to1_xor0 ^ b[3];
  assign arrdiv_fs59_fs_not0 = ~arrdiv_mux2to144_mux2to1_xor0;
  assign arrdiv_fs59_fs_and0 = arrdiv_fs59_fs_not0 & b[3];
  assign arrdiv_fs59_fs_xor1 = arrdiv_fs58_fs_or0 ^ arrdiv_fs59_fs_xor0;
  assign arrdiv_fs59_fs_not1 = ~arrdiv_fs59_fs_xor0;
  assign arrdiv_fs59_fs_and1 = arrdiv_fs59_fs_not1 & arrdiv_fs58_fs_or0;
  assign arrdiv_fs59_fs_or0 = arrdiv_fs59_fs_and1 | arrdiv_fs59_fs_and0;
  assign arrdiv_fs60_fs_xor0 = arrdiv_mux2to145_mux2to1_xor0 ^ b[4];
  assign arrdiv_fs60_fs_not0 = ~arrdiv_mux2to145_mux2to1_xor0;
  assign arrdiv_fs60_fs_and0 = arrdiv_fs60_fs_not0 & b[4];
  assign arrdiv_fs60_fs_xor1 = arrdiv_fs59_fs_or0 ^ arrdiv_fs60_fs_xor0;
  assign arrdiv_fs60_fs_not1 = ~arrdiv_fs60_fs_xor0;
  assign arrdiv_fs60_fs_and1 = arrdiv_fs60_fs_not1 & arrdiv_fs59_fs_or0;
  assign arrdiv_fs60_fs_or0 = arrdiv_fs60_fs_and1 | arrdiv_fs60_fs_and0;
  assign arrdiv_fs61_fs_xor0 = arrdiv_mux2to146_mux2to1_xor0 ^ b[5];
  assign arrdiv_fs61_fs_not0 = ~arrdiv_mux2to146_mux2to1_xor0;
  assign arrdiv_fs61_fs_and0 = arrdiv_fs61_fs_not0 & b[5];
  assign arrdiv_fs61_fs_xor1 = arrdiv_fs60_fs_or0 ^ arrdiv_fs61_fs_xor0;
  assign arrdiv_fs61_fs_not1 = ~arrdiv_fs61_fs_xor0;
  assign arrdiv_fs61_fs_and1 = arrdiv_fs61_fs_not1 & arrdiv_fs60_fs_or0;
  assign arrdiv_fs61_fs_or0 = arrdiv_fs61_fs_and1 | arrdiv_fs61_fs_and0;
  assign arrdiv_fs62_fs_xor0 = arrdiv_mux2to147_mux2to1_xor0 ^ b[6];
  assign arrdiv_fs62_fs_not0 = ~arrdiv_mux2to147_mux2to1_xor0;
  assign arrdiv_fs62_fs_and0 = arrdiv_fs62_fs_not0 & b[6];
  assign arrdiv_fs62_fs_xor1 = arrdiv_fs61_fs_or0 ^ arrdiv_fs62_fs_xor0;
  assign arrdiv_fs62_fs_not1 = ~arrdiv_fs62_fs_xor0;
  assign arrdiv_fs62_fs_and1 = arrdiv_fs62_fs_not1 & arrdiv_fs61_fs_or0;
  assign arrdiv_fs62_fs_or0 = arrdiv_fs62_fs_and1 | arrdiv_fs62_fs_and0;
  assign arrdiv_fs63_fs_xor0 = arrdiv_mux2to148_mux2to1_xor0 ^ b[7];
  assign arrdiv_fs63_fs_not0 = ~arrdiv_mux2to148_mux2to1_xor0;
  assign arrdiv_fs63_fs_and0 = arrdiv_fs63_fs_not0 & b[7];
  assign arrdiv_fs63_fs_xor1 = arrdiv_fs62_fs_or0 ^ arrdiv_fs63_fs_xor0;
  assign arrdiv_fs63_fs_not1 = ~arrdiv_fs63_fs_xor0;
  assign arrdiv_fs63_fs_and1 = arrdiv_fs63_fs_not1 & arrdiv_fs62_fs_or0;
  assign arrdiv_fs63_fs_or0 = arrdiv_fs63_fs_and1 | arrdiv_fs63_fs_and0;
  assign arrdiv_not7 = ~arrdiv_fs63_fs_or0;

  assign arrdiv_out[0] = arrdiv_not7;
  assign arrdiv_out[1] = arrdiv_not6;
  assign arrdiv_out[2] = arrdiv_not5;
  assign arrdiv_out[3] = arrdiv_not4;
  assign arrdiv_out[4] = arrdiv_not3;
  assign arrdiv_out[5] = arrdiv_not2;
  assign arrdiv_out[6] = arrdiv_not1;
  assign arrdiv_out[7] = arrdiv_not0;
endmodule