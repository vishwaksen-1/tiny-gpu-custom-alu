module u_rbs(input [7:0] a, input [7:0] b, output [8:0] u_rbs_out);
  wire u_rbs_hs_hs_xor0;
  wire u_rbs_hs_hs_not0;
  wire u_rbs_hs_hs_xor1;
  wire u_rbs_fs1_fs_xor0;
  wire u_rbs_fs1_fs_not0;
  wire u_rbs_fs1_fs_and0;
  wire u_rbs_fs1_fs_xor1;
  wire u_rbs_fs1_fs_not1;
  wire u_rbs_fs1_fs_and1;
  wire u_rbs_fs1_fs_or0;
  wire u_rbs_fs2_fs_xor0;
  wire u_rbs_fs2_fs_not0;
  wire u_rbs_fs2_fs_and0;
  wire u_rbs_fs2_fs_xor1;
  wire u_rbs_fs2_fs_not1;
  wire u_rbs_fs2_fs_and1;
  wire u_rbs_fs2_fs_or0;
  wire u_rbs_fs3_fs_xor0;
  wire u_rbs_fs3_fs_not0;
  wire u_rbs_fs3_fs_and0;
  wire u_rbs_fs3_fs_xor1;
  wire u_rbs_fs3_fs_not1;
  wire u_rbs_fs3_fs_and1;
  wire u_rbs_fs3_fs_or0;
  wire u_rbs_fs4_fs_xor0;
  wire u_rbs_fs4_fs_not0;
  wire u_rbs_fs4_fs_and0;
  wire u_rbs_fs4_fs_xor1;
  wire u_rbs_fs4_fs_not1;
  wire u_rbs_fs4_fs_and1;
  wire u_rbs_fs4_fs_or0;
  wire u_rbs_fs5_fs_xor0;
  wire u_rbs_fs5_fs_not0;
  wire u_rbs_fs5_fs_and0;
  wire u_rbs_fs5_fs_xor1;
  wire u_rbs_fs5_fs_not1;
  wire u_rbs_fs5_fs_and1;
  wire u_rbs_fs5_fs_or0;
  wire u_rbs_fs6_fs_xor0;
  wire u_rbs_fs6_fs_not0;
  wire u_rbs_fs6_fs_and0;
  wire u_rbs_fs6_fs_xor1;
  wire u_rbs_fs6_fs_not1;
  wire u_rbs_fs6_fs_and1;
  wire u_rbs_fs6_fs_or0;
  wire u_rbs_fs7_fs_xor0;
  wire u_rbs_fs7_fs_not0;
  wire u_rbs_fs7_fs_and0;
  wire u_rbs_fs7_fs_xor1;
  wire u_rbs_fs7_fs_not1;
  wire u_rbs_fs7_fs_and1;
  wire u_rbs_fs7_fs_or0;

  assign u_rbs_hs_hs_xor0 = a[0] ^ b[0];
  assign u_rbs_hs_hs_not0 = ~a[0];
  assign u_rbs_hs_hs_xor1 = u_rbs_hs_hs_not0 & b[0];
  assign u_rbs_fs1_fs_xor0 = a[1] ^ b[1];
  assign u_rbs_fs1_fs_not0 = ~a[1];
  assign u_rbs_fs1_fs_and0 = u_rbs_fs1_fs_not0 & b[1];
  assign u_rbs_fs1_fs_xor1 = u_rbs_hs_hs_xor1 ^ u_rbs_fs1_fs_xor0;
  assign u_rbs_fs1_fs_not1 = ~u_rbs_fs1_fs_xor0;
  assign u_rbs_fs1_fs_and1 = u_rbs_fs1_fs_not1 & u_rbs_hs_hs_xor1;
  assign u_rbs_fs1_fs_or0 = u_rbs_fs1_fs_and1 | u_rbs_fs1_fs_and0;
  assign u_rbs_fs2_fs_xor0 = a[2] ^ b[2];
  assign u_rbs_fs2_fs_not0 = ~a[2];
  assign u_rbs_fs2_fs_and0 = u_rbs_fs2_fs_not0 & b[2];
  assign u_rbs_fs2_fs_xor1 = u_rbs_fs1_fs_or0 ^ u_rbs_fs2_fs_xor0;
  assign u_rbs_fs2_fs_not1 = ~u_rbs_fs2_fs_xor0;
  assign u_rbs_fs2_fs_and1 = u_rbs_fs2_fs_not1 & u_rbs_fs1_fs_or0;
  assign u_rbs_fs2_fs_or0 = u_rbs_fs2_fs_and1 | u_rbs_fs2_fs_and0;
  assign u_rbs_fs3_fs_xor0 = a[3] ^ b[3];
  assign u_rbs_fs3_fs_not0 = ~a[3];
  assign u_rbs_fs3_fs_and0 = u_rbs_fs3_fs_not0 & b[3];
  assign u_rbs_fs3_fs_xor1 = u_rbs_fs2_fs_or0 ^ u_rbs_fs3_fs_xor0;
  assign u_rbs_fs3_fs_not1 = ~u_rbs_fs3_fs_xor0;
  assign u_rbs_fs3_fs_and1 = u_rbs_fs3_fs_not1 & u_rbs_fs2_fs_or0;
  assign u_rbs_fs3_fs_or0 = u_rbs_fs3_fs_and1 | u_rbs_fs3_fs_and0;
  assign u_rbs_fs4_fs_xor0 = a[4] ^ b[4];
  assign u_rbs_fs4_fs_not0 = ~a[4];
  assign u_rbs_fs4_fs_and0 = u_rbs_fs4_fs_not0 & b[4];
  assign u_rbs_fs4_fs_xor1 = u_rbs_fs3_fs_or0 ^ u_rbs_fs4_fs_xor0;
  assign u_rbs_fs4_fs_not1 = ~u_rbs_fs4_fs_xor0;
  assign u_rbs_fs4_fs_and1 = u_rbs_fs4_fs_not1 & u_rbs_fs3_fs_or0;
  assign u_rbs_fs4_fs_or0 = u_rbs_fs4_fs_and1 | u_rbs_fs4_fs_and0;
  assign u_rbs_fs5_fs_xor0 = a[5] ^ b[5];
  assign u_rbs_fs5_fs_not0 = ~a[5];
  assign u_rbs_fs5_fs_and0 = u_rbs_fs5_fs_not0 & b[5];
  assign u_rbs_fs5_fs_xor1 = u_rbs_fs4_fs_or0 ^ u_rbs_fs5_fs_xor0;
  assign u_rbs_fs5_fs_not1 = ~u_rbs_fs5_fs_xor0;
  assign u_rbs_fs5_fs_and1 = u_rbs_fs5_fs_not1 & u_rbs_fs4_fs_or0;
  assign u_rbs_fs5_fs_or0 = u_rbs_fs5_fs_and1 | u_rbs_fs5_fs_and0;
  assign u_rbs_fs6_fs_xor0 = a[6] ^ b[6];
  assign u_rbs_fs6_fs_not0 = ~a[6];
  assign u_rbs_fs6_fs_and0 = u_rbs_fs6_fs_not0 & b[6];
  assign u_rbs_fs6_fs_xor1 = u_rbs_fs5_fs_or0 ^ u_rbs_fs6_fs_xor0;
  assign u_rbs_fs6_fs_not1 = ~u_rbs_fs6_fs_xor0;
  assign u_rbs_fs6_fs_and1 = u_rbs_fs6_fs_not1 & u_rbs_fs5_fs_or0;
  assign u_rbs_fs6_fs_or0 = u_rbs_fs6_fs_and1 | u_rbs_fs6_fs_and0;
  assign u_rbs_fs7_fs_xor0 = a[7] ^ b[7];
  assign u_rbs_fs7_fs_not0 = ~a[7];
  assign u_rbs_fs7_fs_and0 = u_rbs_fs7_fs_not0 & b[7];
  assign u_rbs_fs7_fs_xor1 = u_rbs_fs6_fs_or0 ^ u_rbs_fs7_fs_xor0;
  assign u_rbs_fs7_fs_not1 = ~u_rbs_fs7_fs_xor0;
  assign u_rbs_fs7_fs_and1 = u_rbs_fs7_fs_not1 & u_rbs_fs6_fs_or0;
  assign u_rbs_fs7_fs_or0 = u_rbs_fs7_fs_and1 | u_rbs_fs7_fs_and0;

  assign u_rbs_out[0] = u_rbs_hs_hs_xor0;
  assign u_rbs_out[1] = u_rbs_fs1_fs_xor1;
  assign u_rbs_out[2] = u_rbs_fs2_fs_xor1;
  assign u_rbs_out[3] = u_rbs_fs3_fs_xor1;
  assign u_rbs_out[4] = u_rbs_fs4_fs_xor1;
  assign u_rbs_out[5] = u_rbs_fs5_fs_xor1;
  assign u_rbs_out[6] = u_rbs_fs6_fs_xor1;
  assign u_rbs_out[7] = u_rbs_fs7_fs_xor1;
  assign u_rbs_out[8] = u_rbs_fs7_fs_or0;
endmodule