module u_wallace_cla(input [7:0] a, input [7:0] b, output [15:0] u_wallace_cla_out);
  wire u_wallace_cla_and_0_0;
  wire u_wallace_cla_and_1_0;
  wire u_wallace_cla_and_2_0;
  wire u_wallace_cla_and_3_0;
  wire u_wallace_cla_and_4_0;
  wire u_wallace_cla_and_5_0;
  wire u_wallace_cla_and_6_0;
  wire u_wallace_cla_and_7_0;
  wire u_wallace_cla_and_0_1;
  wire u_wallace_cla_and_1_1;
  wire u_wallace_cla_and_2_1;
  wire u_wallace_cla_and_3_1;
  wire u_wallace_cla_and_4_1;
  wire u_wallace_cla_and_5_1;
  wire u_wallace_cla_and_6_1;
  wire u_wallace_cla_and_7_1;
  wire u_wallace_cla_and_0_2;
  wire u_wallace_cla_and_1_2;
  wire u_wallace_cla_and_2_2;
  wire u_wallace_cla_and_3_2;
  wire u_wallace_cla_and_4_2;
  wire u_wallace_cla_and_5_2;
  wire u_wallace_cla_and_6_2;
  wire u_wallace_cla_and_7_2;
  wire u_wallace_cla_and_0_3;
  wire u_wallace_cla_and_1_3;
  wire u_wallace_cla_and_2_3;
  wire u_wallace_cla_and_3_3;
  wire u_wallace_cla_and_4_3;
  wire u_wallace_cla_and_5_3;
  wire u_wallace_cla_and_6_3;
  wire u_wallace_cla_and_7_3;
  wire u_wallace_cla_and_0_4;
  wire u_wallace_cla_and_1_4;
  wire u_wallace_cla_and_2_4;
  wire u_wallace_cla_and_3_4;
  wire u_wallace_cla_and_4_4;
  wire u_wallace_cla_and_5_4;
  wire u_wallace_cla_and_6_4;
  wire u_wallace_cla_and_7_4;
  wire u_wallace_cla_and_0_5;
  wire u_wallace_cla_and_1_5;
  wire u_wallace_cla_and_2_5;
  wire u_wallace_cla_and_3_5;
  wire u_wallace_cla_and_4_5;
  wire u_wallace_cla_and_5_5;
  wire u_wallace_cla_and_6_5;
  wire u_wallace_cla_and_7_5;
  wire u_wallace_cla_and_0_6;
  wire u_wallace_cla_and_1_6;
  wire u_wallace_cla_and_2_6;
  wire u_wallace_cla_and_3_6;
  wire u_wallace_cla_and_4_6;
  wire u_wallace_cla_and_5_6;
  wire u_wallace_cla_and_6_6;
  wire u_wallace_cla_and_7_6;
  wire u_wallace_cla_and_0_7;
  wire u_wallace_cla_and_1_7;
  wire u_wallace_cla_and_2_7;
  wire u_wallace_cla_and_3_7;
  wire u_wallace_cla_and_4_7;
  wire u_wallace_cla_and_5_7;
  wire u_wallace_cla_and_6_7;
  wire u_wallace_cla_and_7_7;
  wire u_wallace_cla_csa0_csa_component_fa1_fa_xor0;
  wire u_wallace_cla_csa0_csa_component_fa1_fa_and0;
  wire u_wallace_cla_csa0_csa_component_fa2_fa_xor0;
  wire u_wallace_cla_csa0_csa_component_fa2_fa_and0;
  wire u_wallace_cla_csa0_csa_component_fa2_fa_xor1;
  wire u_wallace_cla_csa0_csa_component_fa2_fa_and1;
  wire u_wallace_cla_csa0_csa_component_fa2_fa_or0;
  wire u_wallace_cla_csa0_csa_component_fa3_fa_xor0;
  wire u_wallace_cla_csa0_csa_component_fa3_fa_and0;
  wire u_wallace_cla_csa0_csa_component_fa3_fa_xor1;
  wire u_wallace_cla_csa0_csa_component_fa3_fa_and1;
  wire u_wallace_cla_csa0_csa_component_fa3_fa_or0;
  wire u_wallace_cla_csa0_csa_component_fa4_fa_xor0;
  wire u_wallace_cla_csa0_csa_component_fa4_fa_and0;
  wire u_wallace_cla_csa0_csa_component_fa4_fa_xor1;
  wire u_wallace_cla_csa0_csa_component_fa4_fa_and1;
  wire u_wallace_cla_csa0_csa_component_fa4_fa_or0;
  wire u_wallace_cla_csa0_csa_component_fa5_fa_xor0;
  wire u_wallace_cla_csa0_csa_component_fa5_fa_and0;
  wire u_wallace_cla_csa0_csa_component_fa5_fa_xor1;
  wire u_wallace_cla_csa0_csa_component_fa5_fa_and1;
  wire u_wallace_cla_csa0_csa_component_fa5_fa_or0;
  wire u_wallace_cla_csa0_csa_component_fa6_fa_xor0;
  wire u_wallace_cla_csa0_csa_component_fa6_fa_and0;
  wire u_wallace_cla_csa0_csa_component_fa6_fa_xor1;
  wire u_wallace_cla_csa0_csa_component_fa6_fa_and1;
  wire u_wallace_cla_csa0_csa_component_fa6_fa_or0;
  wire u_wallace_cla_csa0_csa_component_fa7_fa_xor0;
  wire u_wallace_cla_csa0_csa_component_fa7_fa_and0;
  wire u_wallace_cla_csa0_csa_component_fa7_fa_xor1;
  wire u_wallace_cla_csa0_csa_component_fa7_fa_and1;
  wire u_wallace_cla_csa0_csa_component_fa7_fa_or0;
  wire u_wallace_cla_csa0_csa_component_fa8_fa_xor1;
  wire u_wallace_cla_csa0_csa_component_fa8_fa_and1;
  wire u_wallace_cla_csa1_csa_component_fa4_fa_xor0;
  wire u_wallace_cla_csa1_csa_component_fa4_fa_and0;
  wire u_wallace_cla_csa1_csa_component_fa5_fa_xor0;
  wire u_wallace_cla_csa1_csa_component_fa5_fa_and0;
  wire u_wallace_cla_csa1_csa_component_fa5_fa_xor1;
  wire u_wallace_cla_csa1_csa_component_fa5_fa_and1;
  wire u_wallace_cla_csa1_csa_component_fa5_fa_or0;
  wire u_wallace_cla_csa1_csa_component_fa6_fa_xor0;
  wire u_wallace_cla_csa1_csa_component_fa6_fa_and0;
  wire u_wallace_cla_csa1_csa_component_fa6_fa_xor1;
  wire u_wallace_cla_csa1_csa_component_fa6_fa_and1;
  wire u_wallace_cla_csa1_csa_component_fa6_fa_or0;
  wire u_wallace_cla_csa1_csa_component_fa7_fa_xor0;
  wire u_wallace_cla_csa1_csa_component_fa7_fa_and0;
  wire u_wallace_cla_csa1_csa_component_fa7_fa_xor1;
  wire u_wallace_cla_csa1_csa_component_fa7_fa_and1;
  wire u_wallace_cla_csa1_csa_component_fa7_fa_or0;
  wire u_wallace_cla_csa1_csa_component_fa8_fa_xor0;
  wire u_wallace_cla_csa1_csa_component_fa8_fa_and0;
  wire u_wallace_cla_csa1_csa_component_fa8_fa_xor1;
  wire u_wallace_cla_csa1_csa_component_fa8_fa_and1;
  wire u_wallace_cla_csa1_csa_component_fa8_fa_or0;
  wire u_wallace_cla_csa1_csa_component_fa9_fa_xor0;
  wire u_wallace_cla_csa1_csa_component_fa9_fa_and0;
  wire u_wallace_cla_csa1_csa_component_fa9_fa_xor1;
  wire u_wallace_cla_csa1_csa_component_fa9_fa_and1;
  wire u_wallace_cla_csa1_csa_component_fa9_fa_or0;
  wire u_wallace_cla_csa1_csa_component_fa10_fa_xor0;
  wire u_wallace_cla_csa1_csa_component_fa10_fa_and0;
  wire u_wallace_cla_csa1_csa_component_fa10_fa_xor1;
  wire u_wallace_cla_csa1_csa_component_fa10_fa_and1;
  wire u_wallace_cla_csa1_csa_component_fa10_fa_or0;
  wire u_wallace_cla_csa1_csa_component_fa11_fa_xor1;
  wire u_wallace_cla_csa1_csa_component_fa11_fa_and1;
  wire u_wallace_cla_csa2_csa_component_fa2_fa_xor0;
  wire u_wallace_cla_csa2_csa_component_fa2_fa_and0;
  wire u_wallace_cla_csa2_csa_component_fa3_fa_xor0;
  wire u_wallace_cla_csa2_csa_component_fa3_fa_and0;
  wire u_wallace_cla_csa2_csa_component_fa3_fa_xor1;
  wire u_wallace_cla_csa2_csa_component_fa3_fa_and1;
  wire u_wallace_cla_csa2_csa_component_fa3_fa_or0;
  wire u_wallace_cla_csa2_csa_component_fa4_fa_xor0;
  wire u_wallace_cla_csa2_csa_component_fa4_fa_and0;
  wire u_wallace_cla_csa2_csa_component_fa4_fa_xor1;
  wire u_wallace_cla_csa2_csa_component_fa4_fa_and1;
  wire u_wallace_cla_csa2_csa_component_fa4_fa_or0;
  wire u_wallace_cla_csa2_csa_component_fa5_fa_xor0;
  wire u_wallace_cla_csa2_csa_component_fa5_fa_and0;
  wire u_wallace_cla_csa2_csa_component_fa5_fa_xor1;
  wire u_wallace_cla_csa2_csa_component_fa5_fa_and1;
  wire u_wallace_cla_csa2_csa_component_fa5_fa_or0;
  wire u_wallace_cla_csa2_csa_component_fa6_fa_xor0;
  wire u_wallace_cla_csa2_csa_component_fa6_fa_and0;
  wire u_wallace_cla_csa2_csa_component_fa6_fa_xor1;
  wire u_wallace_cla_csa2_csa_component_fa6_fa_and1;
  wire u_wallace_cla_csa2_csa_component_fa6_fa_or0;
  wire u_wallace_cla_csa2_csa_component_fa7_fa_xor0;
  wire u_wallace_cla_csa2_csa_component_fa7_fa_and0;
  wire u_wallace_cla_csa2_csa_component_fa7_fa_xor1;
  wire u_wallace_cla_csa2_csa_component_fa7_fa_and1;
  wire u_wallace_cla_csa2_csa_component_fa7_fa_or0;
  wire u_wallace_cla_csa2_csa_component_fa8_fa_xor0;
  wire u_wallace_cla_csa2_csa_component_fa8_fa_and0;
  wire u_wallace_cla_csa2_csa_component_fa8_fa_xor1;
  wire u_wallace_cla_csa2_csa_component_fa8_fa_and1;
  wire u_wallace_cla_csa2_csa_component_fa8_fa_or0;
  wire u_wallace_cla_csa2_csa_component_fa9_fa_xor0;
  wire u_wallace_cla_csa2_csa_component_fa9_fa_and0;
  wire u_wallace_cla_csa2_csa_component_fa9_fa_xor1;
  wire u_wallace_cla_csa2_csa_component_fa9_fa_and1;
  wire u_wallace_cla_csa2_csa_component_fa9_fa_or0;
  wire u_wallace_cla_csa3_csa_component_fa6_fa_xor0;
  wire u_wallace_cla_csa3_csa_component_fa6_fa_and0;
  wire u_wallace_cla_csa3_csa_component_fa7_fa_xor0;
  wire u_wallace_cla_csa3_csa_component_fa7_fa_and0;
  wire u_wallace_cla_csa3_csa_component_fa7_fa_xor1;
  wire u_wallace_cla_csa3_csa_component_fa7_fa_and1;
  wire u_wallace_cla_csa3_csa_component_fa7_fa_or0;
  wire u_wallace_cla_csa3_csa_component_fa8_fa_xor0;
  wire u_wallace_cla_csa3_csa_component_fa8_fa_and0;
  wire u_wallace_cla_csa3_csa_component_fa8_fa_xor1;
  wire u_wallace_cla_csa3_csa_component_fa8_fa_and1;
  wire u_wallace_cla_csa3_csa_component_fa8_fa_or0;
  wire u_wallace_cla_csa3_csa_component_fa9_fa_xor0;
  wire u_wallace_cla_csa3_csa_component_fa9_fa_and0;
  wire u_wallace_cla_csa3_csa_component_fa9_fa_xor1;
  wire u_wallace_cla_csa3_csa_component_fa9_fa_and1;
  wire u_wallace_cla_csa3_csa_component_fa9_fa_or0;
  wire u_wallace_cla_csa3_csa_component_fa10_fa_xor0;
  wire u_wallace_cla_csa3_csa_component_fa10_fa_and0;
  wire u_wallace_cla_csa3_csa_component_fa10_fa_xor1;
  wire u_wallace_cla_csa3_csa_component_fa10_fa_and1;
  wire u_wallace_cla_csa3_csa_component_fa10_fa_or0;
  wire u_wallace_cla_csa3_csa_component_fa11_fa_xor0;
  wire u_wallace_cla_csa3_csa_component_fa11_fa_and0;
  wire u_wallace_cla_csa3_csa_component_fa11_fa_xor1;
  wire u_wallace_cla_csa3_csa_component_fa11_fa_and1;
  wire u_wallace_cla_csa3_csa_component_fa11_fa_or0;
  wire u_wallace_cla_csa3_csa_component_fa12_fa_xor0;
  wire u_wallace_cla_csa3_csa_component_fa12_fa_and0;
  wire u_wallace_cla_csa3_csa_component_fa12_fa_xor1;
  wire u_wallace_cla_csa3_csa_component_fa12_fa_and1;
  wire u_wallace_cla_csa3_csa_component_fa12_fa_or0;
  wire u_wallace_cla_csa3_csa_component_fa13_fa_xor1;
  wire u_wallace_cla_csa3_csa_component_fa13_fa_and1;
  wire u_wallace_cla_csa4_csa_component_fa3_fa_xor0;
  wire u_wallace_cla_csa4_csa_component_fa3_fa_and0;
  wire u_wallace_cla_csa4_csa_component_fa4_fa_xor0;
  wire u_wallace_cla_csa4_csa_component_fa4_fa_and0;
  wire u_wallace_cla_csa4_csa_component_fa5_fa_xor0;
  wire u_wallace_cla_csa4_csa_component_fa5_fa_and0;
  wire u_wallace_cla_csa4_csa_component_fa5_fa_xor1;
  wire u_wallace_cla_csa4_csa_component_fa5_fa_and1;
  wire u_wallace_cla_csa4_csa_component_fa5_fa_or0;
  wire u_wallace_cla_csa4_csa_component_fa6_fa_xor0;
  wire u_wallace_cla_csa4_csa_component_fa6_fa_and0;
  wire u_wallace_cla_csa4_csa_component_fa6_fa_xor1;
  wire u_wallace_cla_csa4_csa_component_fa6_fa_and1;
  wire u_wallace_cla_csa4_csa_component_fa6_fa_or0;
  wire u_wallace_cla_csa4_csa_component_fa7_fa_xor0;
  wire u_wallace_cla_csa4_csa_component_fa7_fa_and0;
  wire u_wallace_cla_csa4_csa_component_fa7_fa_xor1;
  wire u_wallace_cla_csa4_csa_component_fa7_fa_and1;
  wire u_wallace_cla_csa4_csa_component_fa7_fa_or0;
  wire u_wallace_cla_csa4_csa_component_fa8_fa_xor0;
  wire u_wallace_cla_csa4_csa_component_fa8_fa_and0;
  wire u_wallace_cla_csa4_csa_component_fa8_fa_xor1;
  wire u_wallace_cla_csa4_csa_component_fa8_fa_and1;
  wire u_wallace_cla_csa4_csa_component_fa8_fa_or0;
  wire u_wallace_cla_csa4_csa_component_fa9_fa_xor0;
  wire u_wallace_cla_csa4_csa_component_fa9_fa_and0;
  wire u_wallace_cla_csa4_csa_component_fa9_fa_xor1;
  wire u_wallace_cla_csa4_csa_component_fa9_fa_and1;
  wire u_wallace_cla_csa4_csa_component_fa9_fa_or0;
  wire u_wallace_cla_csa4_csa_component_fa10_fa_xor0;
  wire u_wallace_cla_csa4_csa_component_fa10_fa_and0;
  wire u_wallace_cla_csa4_csa_component_fa10_fa_xor1;
  wire u_wallace_cla_csa4_csa_component_fa10_fa_and1;
  wire u_wallace_cla_csa4_csa_component_fa10_fa_or0;
  wire u_wallace_cla_csa4_csa_component_fa11_fa_xor1;
  wire u_wallace_cla_csa4_csa_component_fa11_fa_and1;
  wire u_wallace_cla_csa4_csa_component_fa12_fa_xor1;
  wire u_wallace_cla_csa4_csa_component_fa12_fa_and1;
  wire u_wallace_cla_csa5_csa_component_fa4_fa_xor0;
  wire u_wallace_cla_csa5_csa_component_fa4_fa_and0;
  wire u_wallace_cla_csa5_csa_component_fa5_fa_xor0;
  wire u_wallace_cla_csa5_csa_component_fa5_fa_and0;
  wire u_wallace_cla_csa5_csa_component_fa6_fa_xor0;
  wire u_wallace_cla_csa5_csa_component_fa6_fa_and0;
  wire u_wallace_cla_csa5_csa_component_fa7_fa_xor0;
  wire u_wallace_cla_csa5_csa_component_fa7_fa_and0;
  wire u_wallace_cla_csa5_csa_component_fa7_fa_xor1;
  wire u_wallace_cla_csa5_csa_component_fa7_fa_and1;
  wire u_wallace_cla_csa5_csa_component_fa7_fa_or0;
  wire u_wallace_cla_csa5_csa_component_fa8_fa_xor0;
  wire u_wallace_cla_csa5_csa_component_fa8_fa_and0;
  wire u_wallace_cla_csa5_csa_component_fa8_fa_xor1;
  wire u_wallace_cla_csa5_csa_component_fa8_fa_and1;
  wire u_wallace_cla_csa5_csa_component_fa8_fa_or0;
  wire u_wallace_cla_csa5_csa_component_fa9_fa_xor0;
  wire u_wallace_cla_csa5_csa_component_fa9_fa_and0;
  wire u_wallace_cla_csa5_csa_component_fa9_fa_xor1;
  wire u_wallace_cla_csa5_csa_component_fa9_fa_and1;
  wire u_wallace_cla_csa5_csa_component_fa9_fa_or0;
  wire u_wallace_cla_csa5_csa_component_fa10_fa_xor0;
  wire u_wallace_cla_csa5_csa_component_fa10_fa_and0;
  wire u_wallace_cla_csa5_csa_component_fa10_fa_xor1;
  wire u_wallace_cla_csa5_csa_component_fa10_fa_and1;
  wire u_wallace_cla_csa5_csa_component_fa10_fa_or0;
  wire u_wallace_cla_csa5_csa_component_fa11_fa_xor0;
  wire u_wallace_cla_csa5_csa_component_fa11_fa_and0;
  wire u_wallace_cla_csa5_csa_component_fa11_fa_xor1;
  wire u_wallace_cla_csa5_csa_component_fa11_fa_and1;
  wire u_wallace_cla_csa5_csa_component_fa11_fa_or0;
  wire u_wallace_cla_csa5_csa_component_fa12_fa_xor0;
  wire u_wallace_cla_csa5_csa_component_fa12_fa_and0;
  wire u_wallace_cla_csa5_csa_component_fa12_fa_xor1;
  wire u_wallace_cla_csa5_csa_component_fa12_fa_and1;
  wire u_wallace_cla_csa5_csa_component_fa12_fa_or0;
  wire u_wallace_cla_csa5_csa_component_fa13_fa_xor0;
  wire u_wallace_cla_csa5_csa_component_fa13_fa_and0;
  wire u_wallace_cla_csa5_csa_component_fa13_fa_xor1;
  wire u_wallace_cla_csa5_csa_component_fa13_fa_and1;
  wire u_wallace_cla_csa5_csa_component_fa13_fa_or0;
  wire u_wallace_cla_csa5_csa_component_fa14_fa_xor1;
  wire u_wallace_cla_csa5_csa_component_fa14_fa_and1;
  wire u_wallace_cla_u_cla16_and0_2_0_1_0;
  wire u_wallace_cla_u_cla16_and0_3_0_1_1;
  wire u_wallace_cla_u_cla16_and0_3_1_1_2;
  wire u_wallace_cla_u_cla16_pg_logic5_pg_logic_or0;
  wire u_wallace_cla_u_cla16_pg_logic5_pg_logic_and0;
  wire u_wallace_cla_u_cla16_pg_logic5_pg_logic_xor0;
  wire u_wallace_cla_u_cla16_pg_logic6_pg_logic_or0;
  wire u_wallace_cla_u_cla16_pg_logic6_pg_logic_and0;
  wire u_wallace_cla_u_cla16_pg_logic6_pg_logic_xor0;
  wire u_wallace_cla_u_cla16_xor6;
  wire u_wallace_cla_u_cla16_and1_2_0_1_3;
  wire u_wallace_cla_u_cla16_and1_2_2_0_4;
  wire u_wallace_cla_u_cla16_or1_2_2_0;
  wire u_wallace_cla_u_cla16_pg_logic7_pg_logic_or0;
  wire u_wallace_cla_u_cla16_pg_logic7_pg_logic_and0;
  wire u_wallace_cla_u_cla16_pg_logic7_pg_logic_xor0;
  wire u_wallace_cla_u_cla16_xor7;
  wire u_wallace_cla_u_cla16_and1_3_0_1_5;
  wire u_wallace_cla_u_cla16_and1_3_1_1_6;
  wire u_wallace_cla_u_cla16_and1_3_2_0_7;
  wire u_wallace_cla_u_cla16_and1_3_2_1_8;
  wire u_wallace_cla_u_cla16_and1_3_3_0_9;
  wire u_wallace_cla_u_cla16_orred1_3_3__2_1;
  wire u_wallace_cla_u_cla16_or1_3_3_2;
  wire u_wallace_cla_u_cla16_pg_logic8_pg_logic_or0;
  wire u_wallace_cla_u_cla16_pg_logic8_pg_logic_and0;
  wire u_wallace_cla_u_cla16_pg_logic8_pg_logic_xor0;
  wire u_wallace_cla_u_cla16_xor8;
  wire u_wallace_cla_u_cla16_and2_0_0_0_10;
  wire u_wallace_cla_u_cla16_or2_0_0_3;
  wire u_wallace_cla_u_cla16_pg_logic9_pg_logic_or0;
  wire u_wallace_cla_u_cla16_pg_logic9_pg_logic_and0;
  wire u_wallace_cla_u_cla16_pg_logic9_pg_logic_xor0;
  wire u_wallace_cla_u_cla16_xor9;
  wire u_wallace_cla_u_cla16_and2_1_0_0_11;
  wire u_wallace_cla_u_cla16_and2_1_0_1_12;
  wire u_wallace_cla_u_cla16_and2_1_1_0_13;
  wire u_wallace_cla_u_cla16_orred2_1_1__0_4;
  wire u_wallace_cla_u_cla16_or2_1_1_5;
  wire u_wallace_cla_u_cla16_pg_logic10_pg_logic_or0;
  wire u_wallace_cla_u_cla16_pg_logic10_pg_logic_and0;
  wire u_wallace_cla_u_cla16_pg_logic10_pg_logic_xor0;
  wire u_wallace_cla_u_cla16_xor10;
  wire u_wallace_cla_u_cla16_and2_2_0_0_14;
  wire u_wallace_cla_u_cla16_and2_2_0_1_15;
  wire u_wallace_cla_u_cla16_and2_2_0_2_16;
  wire u_wallace_cla_u_cla16_and2_2_1_0_17;
  wire u_wallace_cla_u_cla16_and2_2_1_1_18;
  wire u_wallace_cla_u_cla16_and2_2_2_0_19;
  wire u_wallace_cla_u_cla16_orred2_2_2__0_6;
  wire u_wallace_cla_u_cla16_orred2_2_2__1_7;
  wire u_wallace_cla_u_cla16_or2_2_2_8;
  wire u_wallace_cla_u_cla16_pg_logic11_pg_logic_or0;
  wire u_wallace_cla_u_cla16_pg_logic11_pg_logic_and0;
  wire u_wallace_cla_u_cla16_pg_logic11_pg_logic_xor0;
  wire u_wallace_cla_u_cla16_xor11;
  wire u_wallace_cla_u_cla16_and2_3_0_0_20;
  wire u_wallace_cla_u_cla16_and2_3_0_1_21;
  wire u_wallace_cla_u_cla16_and2_3_0_2_22;
  wire u_wallace_cla_u_cla16_and2_3_0_3_23;
  wire u_wallace_cla_u_cla16_and2_3_1_0_24;
  wire u_wallace_cla_u_cla16_and2_3_1_1_25;
  wire u_wallace_cla_u_cla16_and2_3_1_2_26;
  wire u_wallace_cla_u_cla16_and2_3_2_0_27;
  wire u_wallace_cla_u_cla16_and2_3_2_1_28;
  wire u_wallace_cla_u_cla16_and2_3_3_0_29;
  wire u_wallace_cla_u_cla16_orred2_3_3__0_9;
  wire u_wallace_cla_u_cla16_orred2_3_3__1_10;
  wire u_wallace_cla_u_cla16_orred2_3_3__2_11;
  wire u_wallace_cla_u_cla16_or2_3_3_12;
  wire u_wallace_cla_u_cla16_pg_logic12_pg_logic_or0;
  wire u_wallace_cla_u_cla16_pg_logic12_pg_logic_and0;
  wire u_wallace_cla_u_cla16_pg_logic12_pg_logic_xor0;
  wire u_wallace_cla_u_cla16_xor12;
  wire u_wallace_cla_u_cla16_and3_0_0_0_30;
  wire u_wallace_cla_u_cla16_or3_0_0_13;
  wire u_wallace_cla_u_cla16_pg_logic13_pg_logic_or0;
  wire u_wallace_cla_u_cla16_pg_logic13_pg_logic_and0;
  wire u_wallace_cla_u_cla16_pg_logic13_pg_logic_xor0;
  wire u_wallace_cla_u_cla16_xor13;
  wire u_wallace_cla_u_cla16_and3_1_0_0_31;
  wire u_wallace_cla_u_cla16_and3_1_0_1_32;
  wire u_wallace_cla_u_cla16_and3_1_1_0_33;
  wire u_wallace_cla_u_cla16_orred3_1_1__0_14;
  wire u_wallace_cla_u_cla16_or3_1_1_15;
  wire u_wallace_cla_u_cla16_pg_logic14_pg_logic_or0;
  wire u_wallace_cla_u_cla16_pg_logic14_pg_logic_and0;
  wire u_wallace_cla_u_cla16_pg_logic14_pg_logic_xor0;
  wire u_wallace_cla_u_cla16_xor14;
  wire u_wallace_cla_u_cla16_and3_2_0_0_34;
  wire u_wallace_cla_u_cla16_and3_2_0_1_35;
  wire u_wallace_cla_u_cla16_and3_2_0_2_36;
  wire u_wallace_cla_u_cla16_and3_2_1_0_37;
  wire u_wallace_cla_u_cla16_and3_2_1_1_38;
  wire u_wallace_cla_u_cla16_and3_2_2_0_39;
  wire u_wallace_cla_u_cla16_orred3_2_2__0_16;
  wire u_wallace_cla_u_cla16_orred3_2_2__1_17;
  wire u_wallace_cla_u_cla16_or3_2_2_18;
  wire u_wallace_cla_u_cla16_xor15;
  wire u_wallace_cla_u_cla16_and3_3_0_0_40;
  wire u_wallace_cla_u_cla16_and3_3_0_1_41;
  wire u_wallace_cla_u_cla16_and3_3_0_2_42;
  wire u_wallace_cla_u_cla16_and3_3_0_3_43;
  wire u_wallace_cla_u_cla16_and3_3_1_0_44;
  wire u_wallace_cla_u_cla16_and3_3_1_1_45;
  wire u_wallace_cla_u_cla16_and3_3_1_2_46;
  wire u_wallace_cla_u_cla16_and3_3_2_0_47;
  wire u_wallace_cla_u_cla16_and3_3_2_1_48;
  wire u_wallace_cla_u_cla16_and3_3_3_0_49;
  wire u_wallace_cla_u_cla16_orred3_3_3__0_19;
  wire u_wallace_cla_u_cla16_orred3_3_3__1_20;
  wire u_wallace_cla_u_cla16_orred3_3_3__2_21;

  assign u_wallace_cla_and_0_0 = a[0] & b[0];
  assign u_wallace_cla_and_1_0 = a[1] & b[0];
  assign u_wallace_cla_and_2_0 = a[2] & b[0];
  assign u_wallace_cla_and_3_0 = a[3] & b[0];
  assign u_wallace_cla_and_4_0 = a[4] & b[0];
  assign u_wallace_cla_and_5_0 = a[5] & b[0];
  assign u_wallace_cla_and_6_0 = a[6] & b[0];
  assign u_wallace_cla_and_7_0 = a[7] & b[0];
  assign u_wallace_cla_and_0_1 = a[0] & b[1];
  assign u_wallace_cla_and_1_1 = a[1] & b[1];
  assign u_wallace_cla_and_2_1 = a[2] & b[1];
  assign u_wallace_cla_and_3_1 = a[3] & b[1];
  assign u_wallace_cla_and_4_1 = a[4] & b[1];
  assign u_wallace_cla_and_5_1 = a[5] & b[1];
  assign u_wallace_cla_and_6_1 = a[6] & b[1];
  assign u_wallace_cla_and_7_1 = a[7] & b[1];
  assign u_wallace_cla_and_0_2 = a[0] & b[2];
  assign u_wallace_cla_and_1_2 = a[1] & b[2];
  assign u_wallace_cla_and_2_2 = a[2] & b[2];
  assign u_wallace_cla_and_3_2 = a[3] & b[2];
  assign u_wallace_cla_and_4_2 = a[4] & b[2];
  assign u_wallace_cla_and_5_2 = a[5] & b[2];
  assign u_wallace_cla_and_6_2 = a[6] & b[2];
  assign u_wallace_cla_and_7_2 = a[7] & b[2];
  assign u_wallace_cla_and_0_3 = a[0] & b[3];
  assign u_wallace_cla_and_1_3 = a[1] & b[3];
  assign u_wallace_cla_and_2_3 = a[2] & b[3];
  assign u_wallace_cla_and_3_3 = a[3] & b[3];
  assign u_wallace_cla_and_4_3 = a[4] & b[3];
  assign u_wallace_cla_and_5_3 = a[5] & b[3];
  assign u_wallace_cla_and_6_3 = a[6] & b[3];
  assign u_wallace_cla_and_7_3 = a[7] & b[3];
  assign u_wallace_cla_and_0_4 = a[0] & b[4];
  assign u_wallace_cla_and_1_4 = a[1] & b[4];
  assign u_wallace_cla_and_2_4 = a[2] & b[4];
  assign u_wallace_cla_and_3_4 = a[3] & b[4];
  assign u_wallace_cla_and_4_4 = a[4] & b[4];
  assign u_wallace_cla_and_5_4 = a[5] & b[4];
  assign u_wallace_cla_and_6_4 = a[6] & b[4];
  assign u_wallace_cla_and_7_4 = a[7] & b[4];
  assign u_wallace_cla_and_0_5 = a[0] & b[5];
  assign u_wallace_cla_and_1_5 = a[1] & b[5];
  assign u_wallace_cla_and_2_5 = a[2] & b[5];
  assign u_wallace_cla_and_3_5 = a[3] & b[5];
  assign u_wallace_cla_and_4_5 = a[4] & b[5];
  assign u_wallace_cla_and_5_5 = a[5] & b[5];
  assign u_wallace_cla_and_6_5 = a[6] & b[5];
  assign u_wallace_cla_and_7_5 = a[7] & b[5];
  assign u_wallace_cla_and_0_6 = a[0] & b[6];
  assign u_wallace_cla_and_1_6 = a[1] & b[6];
  assign u_wallace_cla_and_2_6 = a[2] & b[6];
  assign u_wallace_cla_and_3_6 = a[3] & b[6];
  assign u_wallace_cla_and_4_6 = a[4] & b[6];
  assign u_wallace_cla_and_5_6 = a[5] & b[6];
  assign u_wallace_cla_and_6_6 = a[6] & b[6];
  assign u_wallace_cla_and_7_6 = a[7] & b[6];
  assign u_wallace_cla_and_0_7 = a[0] & b[7];
  assign u_wallace_cla_and_1_7 = a[1] & b[7];
  assign u_wallace_cla_and_2_7 = a[2] & b[7];
  assign u_wallace_cla_and_3_7 = a[3] & b[7];
  assign u_wallace_cla_and_4_7 = a[4] & b[7];
  assign u_wallace_cla_and_5_7 = a[5] & b[7];
  assign u_wallace_cla_and_6_7 = a[6] & b[7];
  assign u_wallace_cla_and_7_7 = a[7] & b[7];
  assign u_wallace_cla_csa0_csa_component_fa1_fa_xor0 = u_wallace_cla_and_1_0 ^ u_wallace_cla_and_0_1;
  assign u_wallace_cla_csa0_csa_component_fa1_fa_and0 = u_wallace_cla_and_1_0 & u_wallace_cla_and_0_1;
  assign u_wallace_cla_csa0_csa_component_fa2_fa_xor0 = u_wallace_cla_and_2_0 ^ u_wallace_cla_and_1_1;
  assign u_wallace_cla_csa0_csa_component_fa2_fa_and0 = u_wallace_cla_and_2_0 & u_wallace_cla_and_1_1;
  assign u_wallace_cla_csa0_csa_component_fa2_fa_xor1 = u_wallace_cla_csa0_csa_component_fa2_fa_xor0 ^ u_wallace_cla_and_0_2;
  assign u_wallace_cla_csa0_csa_component_fa2_fa_and1 = u_wallace_cla_csa0_csa_component_fa2_fa_xor0 & u_wallace_cla_and_0_2;
  assign u_wallace_cla_csa0_csa_component_fa2_fa_or0 = u_wallace_cla_csa0_csa_component_fa2_fa_and0 | u_wallace_cla_csa0_csa_component_fa2_fa_and1;
  assign u_wallace_cla_csa0_csa_component_fa3_fa_xor0 = u_wallace_cla_and_3_0 ^ u_wallace_cla_and_2_1;
  assign u_wallace_cla_csa0_csa_component_fa3_fa_and0 = u_wallace_cla_and_3_0 & u_wallace_cla_and_2_1;
  assign u_wallace_cla_csa0_csa_component_fa3_fa_xor1 = u_wallace_cla_csa0_csa_component_fa3_fa_xor0 ^ u_wallace_cla_and_1_2;
  assign u_wallace_cla_csa0_csa_component_fa3_fa_and1 = u_wallace_cla_csa0_csa_component_fa3_fa_xor0 & u_wallace_cla_and_1_2;
  assign u_wallace_cla_csa0_csa_component_fa3_fa_or0 = u_wallace_cla_csa0_csa_component_fa3_fa_and0 | u_wallace_cla_csa0_csa_component_fa3_fa_and1;
  assign u_wallace_cla_csa0_csa_component_fa4_fa_xor0 = u_wallace_cla_and_4_0 ^ u_wallace_cla_and_3_1;
  assign u_wallace_cla_csa0_csa_component_fa4_fa_and0 = u_wallace_cla_and_4_0 & u_wallace_cla_and_3_1;
  assign u_wallace_cla_csa0_csa_component_fa4_fa_xor1 = u_wallace_cla_csa0_csa_component_fa4_fa_xor0 ^ u_wallace_cla_and_2_2;
  assign u_wallace_cla_csa0_csa_component_fa4_fa_and1 = u_wallace_cla_csa0_csa_component_fa4_fa_xor0 & u_wallace_cla_and_2_2;
  assign u_wallace_cla_csa0_csa_component_fa4_fa_or0 = u_wallace_cla_csa0_csa_component_fa4_fa_and0 | u_wallace_cla_csa0_csa_component_fa4_fa_and1;
  assign u_wallace_cla_csa0_csa_component_fa5_fa_xor0 = u_wallace_cla_and_5_0 ^ u_wallace_cla_and_4_1;
  assign u_wallace_cla_csa0_csa_component_fa5_fa_and0 = u_wallace_cla_and_5_0 & u_wallace_cla_and_4_1;
  assign u_wallace_cla_csa0_csa_component_fa5_fa_xor1 = u_wallace_cla_csa0_csa_component_fa5_fa_xor0 ^ u_wallace_cla_and_3_2;
  assign u_wallace_cla_csa0_csa_component_fa5_fa_and1 = u_wallace_cla_csa0_csa_component_fa5_fa_xor0 & u_wallace_cla_and_3_2;
  assign u_wallace_cla_csa0_csa_component_fa5_fa_or0 = u_wallace_cla_csa0_csa_component_fa5_fa_and0 | u_wallace_cla_csa0_csa_component_fa5_fa_and1;
  assign u_wallace_cla_csa0_csa_component_fa6_fa_xor0 = u_wallace_cla_and_6_0 ^ u_wallace_cla_and_5_1;
  assign u_wallace_cla_csa0_csa_component_fa6_fa_and0 = u_wallace_cla_and_6_0 & u_wallace_cla_and_5_1;
  assign u_wallace_cla_csa0_csa_component_fa6_fa_xor1 = u_wallace_cla_csa0_csa_component_fa6_fa_xor0 ^ u_wallace_cla_and_4_2;
  assign u_wallace_cla_csa0_csa_component_fa6_fa_and1 = u_wallace_cla_csa0_csa_component_fa6_fa_xor0 & u_wallace_cla_and_4_2;
  assign u_wallace_cla_csa0_csa_component_fa6_fa_or0 = u_wallace_cla_csa0_csa_component_fa6_fa_and0 | u_wallace_cla_csa0_csa_component_fa6_fa_and1;
  assign u_wallace_cla_csa0_csa_component_fa7_fa_xor0 = u_wallace_cla_and_7_0 ^ u_wallace_cla_and_6_1;
  assign u_wallace_cla_csa0_csa_component_fa7_fa_and0 = u_wallace_cla_and_7_0 & u_wallace_cla_and_6_1;
  assign u_wallace_cla_csa0_csa_component_fa7_fa_xor1 = u_wallace_cla_csa0_csa_component_fa7_fa_xor0 ^ u_wallace_cla_and_5_2;
  assign u_wallace_cla_csa0_csa_component_fa7_fa_and1 = u_wallace_cla_csa0_csa_component_fa7_fa_xor0 & u_wallace_cla_and_5_2;
  assign u_wallace_cla_csa0_csa_component_fa7_fa_or0 = u_wallace_cla_csa0_csa_component_fa7_fa_and0 | u_wallace_cla_csa0_csa_component_fa7_fa_and1;
  assign u_wallace_cla_csa0_csa_component_fa8_fa_xor1 = u_wallace_cla_and_7_1 ^ u_wallace_cla_and_6_2;
  assign u_wallace_cla_csa0_csa_component_fa8_fa_and1 = u_wallace_cla_and_7_1 & u_wallace_cla_and_6_2;
  assign u_wallace_cla_csa1_csa_component_fa4_fa_xor0 = u_wallace_cla_and_1_3 ^ u_wallace_cla_and_0_4;
  assign u_wallace_cla_csa1_csa_component_fa4_fa_and0 = u_wallace_cla_and_1_3 & u_wallace_cla_and_0_4;
  assign u_wallace_cla_csa1_csa_component_fa5_fa_xor0 = u_wallace_cla_and_2_3 ^ u_wallace_cla_and_1_4;
  assign u_wallace_cla_csa1_csa_component_fa5_fa_and0 = u_wallace_cla_and_2_3 & u_wallace_cla_and_1_4;
  assign u_wallace_cla_csa1_csa_component_fa5_fa_xor1 = u_wallace_cla_csa1_csa_component_fa5_fa_xor0 ^ u_wallace_cla_and_0_5;
  assign u_wallace_cla_csa1_csa_component_fa5_fa_and1 = u_wallace_cla_csa1_csa_component_fa5_fa_xor0 & u_wallace_cla_and_0_5;
  assign u_wallace_cla_csa1_csa_component_fa5_fa_or0 = u_wallace_cla_csa1_csa_component_fa5_fa_and0 | u_wallace_cla_csa1_csa_component_fa5_fa_and1;
  assign u_wallace_cla_csa1_csa_component_fa6_fa_xor0 = u_wallace_cla_and_3_3 ^ u_wallace_cla_and_2_4;
  assign u_wallace_cla_csa1_csa_component_fa6_fa_and0 = u_wallace_cla_and_3_3 & u_wallace_cla_and_2_4;
  assign u_wallace_cla_csa1_csa_component_fa6_fa_xor1 = u_wallace_cla_csa1_csa_component_fa6_fa_xor0 ^ u_wallace_cla_and_1_5;
  assign u_wallace_cla_csa1_csa_component_fa6_fa_and1 = u_wallace_cla_csa1_csa_component_fa6_fa_xor0 & u_wallace_cla_and_1_5;
  assign u_wallace_cla_csa1_csa_component_fa6_fa_or0 = u_wallace_cla_csa1_csa_component_fa6_fa_and0 | u_wallace_cla_csa1_csa_component_fa6_fa_and1;
  assign u_wallace_cla_csa1_csa_component_fa7_fa_xor0 = u_wallace_cla_and_4_3 ^ u_wallace_cla_and_3_4;
  assign u_wallace_cla_csa1_csa_component_fa7_fa_and0 = u_wallace_cla_and_4_3 & u_wallace_cla_and_3_4;
  assign u_wallace_cla_csa1_csa_component_fa7_fa_xor1 = u_wallace_cla_csa1_csa_component_fa7_fa_xor0 ^ u_wallace_cla_and_2_5;
  assign u_wallace_cla_csa1_csa_component_fa7_fa_and1 = u_wallace_cla_csa1_csa_component_fa7_fa_xor0 & u_wallace_cla_and_2_5;
  assign u_wallace_cla_csa1_csa_component_fa7_fa_or0 = u_wallace_cla_csa1_csa_component_fa7_fa_and0 | u_wallace_cla_csa1_csa_component_fa7_fa_and1;
  assign u_wallace_cla_csa1_csa_component_fa8_fa_xor0 = u_wallace_cla_and_5_3 ^ u_wallace_cla_and_4_4;
  assign u_wallace_cla_csa1_csa_component_fa8_fa_and0 = u_wallace_cla_and_5_3 & u_wallace_cla_and_4_4;
  assign u_wallace_cla_csa1_csa_component_fa8_fa_xor1 = u_wallace_cla_csa1_csa_component_fa8_fa_xor0 ^ u_wallace_cla_and_3_5;
  assign u_wallace_cla_csa1_csa_component_fa8_fa_and1 = u_wallace_cla_csa1_csa_component_fa8_fa_xor0 & u_wallace_cla_and_3_5;
  assign u_wallace_cla_csa1_csa_component_fa8_fa_or0 = u_wallace_cla_csa1_csa_component_fa8_fa_and0 | u_wallace_cla_csa1_csa_component_fa8_fa_and1;
  assign u_wallace_cla_csa1_csa_component_fa9_fa_xor0 = u_wallace_cla_and_6_3 ^ u_wallace_cla_and_5_4;
  assign u_wallace_cla_csa1_csa_component_fa9_fa_and0 = u_wallace_cla_and_6_3 & u_wallace_cla_and_5_4;
  assign u_wallace_cla_csa1_csa_component_fa9_fa_xor1 = u_wallace_cla_csa1_csa_component_fa9_fa_xor0 ^ u_wallace_cla_and_4_5;
  assign u_wallace_cla_csa1_csa_component_fa9_fa_and1 = u_wallace_cla_csa1_csa_component_fa9_fa_xor0 & u_wallace_cla_and_4_5;
  assign u_wallace_cla_csa1_csa_component_fa9_fa_or0 = u_wallace_cla_csa1_csa_component_fa9_fa_and0 | u_wallace_cla_csa1_csa_component_fa9_fa_and1;
  assign u_wallace_cla_csa1_csa_component_fa10_fa_xor0 = u_wallace_cla_and_7_3 ^ u_wallace_cla_and_6_4;
  assign u_wallace_cla_csa1_csa_component_fa10_fa_and0 = u_wallace_cla_and_7_3 & u_wallace_cla_and_6_4;
  assign u_wallace_cla_csa1_csa_component_fa10_fa_xor1 = u_wallace_cla_csa1_csa_component_fa10_fa_xor0 ^ u_wallace_cla_and_5_5;
  assign u_wallace_cla_csa1_csa_component_fa10_fa_and1 = u_wallace_cla_csa1_csa_component_fa10_fa_xor0 & u_wallace_cla_and_5_5;
  assign u_wallace_cla_csa1_csa_component_fa10_fa_or0 = u_wallace_cla_csa1_csa_component_fa10_fa_and0 | u_wallace_cla_csa1_csa_component_fa10_fa_and1;
  assign u_wallace_cla_csa1_csa_component_fa11_fa_xor1 = u_wallace_cla_and_7_4 ^ u_wallace_cla_and_6_5;
  assign u_wallace_cla_csa1_csa_component_fa11_fa_and1 = u_wallace_cla_and_7_4 & u_wallace_cla_and_6_5;
  assign u_wallace_cla_csa2_csa_component_fa2_fa_xor0 = u_wallace_cla_csa0_csa_component_fa2_fa_xor1 ^ u_wallace_cla_csa0_csa_component_fa1_fa_and0;
  assign u_wallace_cla_csa2_csa_component_fa2_fa_and0 = u_wallace_cla_csa0_csa_component_fa2_fa_xor1 & u_wallace_cla_csa0_csa_component_fa1_fa_and0;
  assign u_wallace_cla_csa2_csa_component_fa3_fa_xor0 = u_wallace_cla_csa0_csa_component_fa3_fa_xor1 ^ u_wallace_cla_csa0_csa_component_fa2_fa_or0;
  assign u_wallace_cla_csa2_csa_component_fa3_fa_and0 = u_wallace_cla_csa0_csa_component_fa3_fa_xor1 & u_wallace_cla_csa0_csa_component_fa2_fa_or0;
  assign u_wallace_cla_csa2_csa_component_fa3_fa_xor1 = u_wallace_cla_csa2_csa_component_fa3_fa_xor0 ^ u_wallace_cla_and_0_3;
  assign u_wallace_cla_csa2_csa_component_fa3_fa_and1 = u_wallace_cla_csa2_csa_component_fa3_fa_xor0 & u_wallace_cla_and_0_3;
  assign u_wallace_cla_csa2_csa_component_fa3_fa_or0 = u_wallace_cla_csa2_csa_component_fa3_fa_and0 | u_wallace_cla_csa2_csa_component_fa3_fa_and1;
  assign u_wallace_cla_csa2_csa_component_fa4_fa_xor0 = u_wallace_cla_csa0_csa_component_fa4_fa_xor1 ^ u_wallace_cla_csa0_csa_component_fa3_fa_or0;
  assign u_wallace_cla_csa2_csa_component_fa4_fa_and0 = u_wallace_cla_csa0_csa_component_fa4_fa_xor1 & u_wallace_cla_csa0_csa_component_fa3_fa_or0;
  assign u_wallace_cla_csa2_csa_component_fa4_fa_xor1 = u_wallace_cla_csa2_csa_component_fa4_fa_xor0 ^ u_wallace_cla_csa1_csa_component_fa4_fa_xor0;
  assign u_wallace_cla_csa2_csa_component_fa4_fa_and1 = u_wallace_cla_csa2_csa_component_fa4_fa_xor0 & u_wallace_cla_csa1_csa_component_fa4_fa_xor0;
  assign u_wallace_cla_csa2_csa_component_fa4_fa_or0 = u_wallace_cla_csa2_csa_component_fa4_fa_and0 | u_wallace_cla_csa2_csa_component_fa4_fa_and1;
  assign u_wallace_cla_csa2_csa_component_fa5_fa_xor0 = u_wallace_cla_csa0_csa_component_fa5_fa_xor1 ^ u_wallace_cla_csa0_csa_component_fa4_fa_or0;
  assign u_wallace_cla_csa2_csa_component_fa5_fa_and0 = u_wallace_cla_csa0_csa_component_fa5_fa_xor1 & u_wallace_cla_csa0_csa_component_fa4_fa_or0;
  assign u_wallace_cla_csa2_csa_component_fa5_fa_xor1 = u_wallace_cla_csa2_csa_component_fa5_fa_xor0 ^ u_wallace_cla_csa1_csa_component_fa5_fa_xor1;
  assign u_wallace_cla_csa2_csa_component_fa5_fa_and1 = u_wallace_cla_csa2_csa_component_fa5_fa_xor0 & u_wallace_cla_csa1_csa_component_fa5_fa_xor1;
  assign u_wallace_cla_csa2_csa_component_fa5_fa_or0 = u_wallace_cla_csa2_csa_component_fa5_fa_and0 | u_wallace_cla_csa2_csa_component_fa5_fa_and1;
  assign u_wallace_cla_csa2_csa_component_fa6_fa_xor0 = u_wallace_cla_csa0_csa_component_fa6_fa_xor1 ^ u_wallace_cla_csa0_csa_component_fa5_fa_or0;
  assign u_wallace_cla_csa2_csa_component_fa6_fa_and0 = u_wallace_cla_csa0_csa_component_fa6_fa_xor1 & u_wallace_cla_csa0_csa_component_fa5_fa_or0;
  assign u_wallace_cla_csa2_csa_component_fa6_fa_xor1 = u_wallace_cla_csa2_csa_component_fa6_fa_xor0 ^ u_wallace_cla_csa1_csa_component_fa6_fa_xor1;
  assign u_wallace_cla_csa2_csa_component_fa6_fa_and1 = u_wallace_cla_csa2_csa_component_fa6_fa_xor0 & u_wallace_cla_csa1_csa_component_fa6_fa_xor1;
  assign u_wallace_cla_csa2_csa_component_fa6_fa_or0 = u_wallace_cla_csa2_csa_component_fa6_fa_and0 | u_wallace_cla_csa2_csa_component_fa6_fa_and1;
  assign u_wallace_cla_csa2_csa_component_fa7_fa_xor0 = u_wallace_cla_csa0_csa_component_fa7_fa_xor1 ^ u_wallace_cla_csa0_csa_component_fa6_fa_or0;
  assign u_wallace_cla_csa2_csa_component_fa7_fa_and0 = u_wallace_cla_csa0_csa_component_fa7_fa_xor1 & u_wallace_cla_csa0_csa_component_fa6_fa_or0;
  assign u_wallace_cla_csa2_csa_component_fa7_fa_xor1 = u_wallace_cla_csa2_csa_component_fa7_fa_xor0 ^ u_wallace_cla_csa1_csa_component_fa7_fa_xor1;
  assign u_wallace_cla_csa2_csa_component_fa7_fa_and1 = u_wallace_cla_csa2_csa_component_fa7_fa_xor0 & u_wallace_cla_csa1_csa_component_fa7_fa_xor1;
  assign u_wallace_cla_csa2_csa_component_fa7_fa_or0 = u_wallace_cla_csa2_csa_component_fa7_fa_and0 | u_wallace_cla_csa2_csa_component_fa7_fa_and1;
  assign u_wallace_cla_csa2_csa_component_fa8_fa_xor0 = u_wallace_cla_csa0_csa_component_fa8_fa_xor1 ^ u_wallace_cla_csa0_csa_component_fa7_fa_or0;
  assign u_wallace_cla_csa2_csa_component_fa8_fa_and0 = u_wallace_cla_csa0_csa_component_fa8_fa_xor1 & u_wallace_cla_csa0_csa_component_fa7_fa_or0;
  assign u_wallace_cla_csa2_csa_component_fa8_fa_xor1 = u_wallace_cla_csa2_csa_component_fa8_fa_xor0 ^ u_wallace_cla_csa1_csa_component_fa8_fa_xor1;
  assign u_wallace_cla_csa2_csa_component_fa8_fa_and1 = u_wallace_cla_csa2_csa_component_fa8_fa_xor0 & u_wallace_cla_csa1_csa_component_fa8_fa_xor1;
  assign u_wallace_cla_csa2_csa_component_fa8_fa_or0 = u_wallace_cla_csa2_csa_component_fa8_fa_and0 | u_wallace_cla_csa2_csa_component_fa8_fa_and1;
  assign u_wallace_cla_csa2_csa_component_fa9_fa_xor0 = u_wallace_cla_and_7_2 ^ u_wallace_cla_csa0_csa_component_fa8_fa_and1;
  assign u_wallace_cla_csa2_csa_component_fa9_fa_and0 = u_wallace_cla_and_7_2 & u_wallace_cla_csa0_csa_component_fa8_fa_and1;
  assign u_wallace_cla_csa2_csa_component_fa9_fa_xor1 = u_wallace_cla_csa2_csa_component_fa9_fa_xor0 ^ u_wallace_cla_csa1_csa_component_fa9_fa_xor1;
  assign u_wallace_cla_csa2_csa_component_fa9_fa_and1 = u_wallace_cla_csa2_csa_component_fa9_fa_xor0 & u_wallace_cla_csa1_csa_component_fa9_fa_xor1;
  assign u_wallace_cla_csa2_csa_component_fa9_fa_or0 = u_wallace_cla_csa2_csa_component_fa9_fa_and0 | u_wallace_cla_csa2_csa_component_fa9_fa_and1;
  assign u_wallace_cla_csa3_csa_component_fa6_fa_xor0 = u_wallace_cla_csa1_csa_component_fa5_fa_or0 ^ u_wallace_cla_and_0_6;
  assign u_wallace_cla_csa3_csa_component_fa6_fa_and0 = u_wallace_cla_csa1_csa_component_fa5_fa_or0 & u_wallace_cla_and_0_6;
  assign u_wallace_cla_csa3_csa_component_fa7_fa_xor0 = u_wallace_cla_csa1_csa_component_fa6_fa_or0 ^ u_wallace_cla_and_1_6;
  assign u_wallace_cla_csa3_csa_component_fa7_fa_and0 = u_wallace_cla_csa1_csa_component_fa6_fa_or0 & u_wallace_cla_and_1_6;
  assign u_wallace_cla_csa3_csa_component_fa7_fa_xor1 = u_wallace_cla_csa3_csa_component_fa7_fa_xor0 ^ u_wallace_cla_and_0_7;
  assign u_wallace_cla_csa3_csa_component_fa7_fa_and1 = u_wallace_cla_csa3_csa_component_fa7_fa_xor0 & u_wallace_cla_and_0_7;
  assign u_wallace_cla_csa3_csa_component_fa7_fa_or0 = u_wallace_cla_csa3_csa_component_fa7_fa_and0 | u_wallace_cla_csa3_csa_component_fa7_fa_and1;
  assign u_wallace_cla_csa3_csa_component_fa8_fa_xor0 = u_wallace_cla_csa1_csa_component_fa7_fa_or0 ^ u_wallace_cla_and_2_6;
  assign u_wallace_cla_csa3_csa_component_fa8_fa_and0 = u_wallace_cla_csa1_csa_component_fa7_fa_or0 & u_wallace_cla_and_2_6;
  assign u_wallace_cla_csa3_csa_component_fa8_fa_xor1 = u_wallace_cla_csa3_csa_component_fa8_fa_xor0 ^ u_wallace_cla_and_1_7;
  assign u_wallace_cla_csa3_csa_component_fa8_fa_and1 = u_wallace_cla_csa3_csa_component_fa8_fa_xor0 & u_wallace_cla_and_1_7;
  assign u_wallace_cla_csa3_csa_component_fa8_fa_or0 = u_wallace_cla_csa3_csa_component_fa8_fa_and0 | u_wallace_cla_csa3_csa_component_fa8_fa_and1;
  assign u_wallace_cla_csa3_csa_component_fa9_fa_xor0 = u_wallace_cla_csa1_csa_component_fa8_fa_or0 ^ u_wallace_cla_and_3_6;
  assign u_wallace_cla_csa3_csa_component_fa9_fa_and0 = u_wallace_cla_csa1_csa_component_fa8_fa_or0 & u_wallace_cla_and_3_6;
  assign u_wallace_cla_csa3_csa_component_fa9_fa_xor1 = u_wallace_cla_csa3_csa_component_fa9_fa_xor0 ^ u_wallace_cla_and_2_7;
  assign u_wallace_cla_csa3_csa_component_fa9_fa_and1 = u_wallace_cla_csa3_csa_component_fa9_fa_xor0 & u_wallace_cla_and_2_7;
  assign u_wallace_cla_csa3_csa_component_fa9_fa_or0 = u_wallace_cla_csa3_csa_component_fa9_fa_and0 | u_wallace_cla_csa3_csa_component_fa9_fa_and1;
  assign u_wallace_cla_csa3_csa_component_fa10_fa_xor0 = u_wallace_cla_csa1_csa_component_fa9_fa_or0 ^ u_wallace_cla_and_4_6;
  assign u_wallace_cla_csa3_csa_component_fa10_fa_and0 = u_wallace_cla_csa1_csa_component_fa9_fa_or0 & u_wallace_cla_and_4_6;
  assign u_wallace_cla_csa3_csa_component_fa10_fa_xor1 = u_wallace_cla_csa3_csa_component_fa10_fa_xor0 ^ u_wallace_cla_and_3_7;
  assign u_wallace_cla_csa3_csa_component_fa10_fa_and1 = u_wallace_cla_csa3_csa_component_fa10_fa_xor0 & u_wallace_cla_and_3_7;
  assign u_wallace_cla_csa3_csa_component_fa10_fa_or0 = u_wallace_cla_csa3_csa_component_fa10_fa_and0 | u_wallace_cla_csa3_csa_component_fa10_fa_and1;
  assign u_wallace_cla_csa3_csa_component_fa11_fa_xor0 = u_wallace_cla_csa1_csa_component_fa10_fa_or0 ^ u_wallace_cla_and_5_6;
  assign u_wallace_cla_csa3_csa_component_fa11_fa_and0 = u_wallace_cla_csa1_csa_component_fa10_fa_or0 & u_wallace_cla_and_5_6;
  assign u_wallace_cla_csa3_csa_component_fa11_fa_xor1 = u_wallace_cla_csa3_csa_component_fa11_fa_xor0 ^ u_wallace_cla_and_4_7;
  assign u_wallace_cla_csa3_csa_component_fa11_fa_and1 = u_wallace_cla_csa3_csa_component_fa11_fa_xor0 & u_wallace_cla_and_4_7;
  assign u_wallace_cla_csa3_csa_component_fa11_fa_or0 = u_wallace_cla_csa3_csa_component_fa11_fa_and0 | u_wallace_cla_csa3_csa_component_fa11_fa_and1;
  assign u_wallace_cla_csa3_csa_component_fa12_fa_xor0 = u_wallace_cla_csa1_csa_component_fa11_fa_and1 ^ u_wallace_cla_and_6_6;
  assign u_wallace_cla_csa3_csa_component_fa12_fa_and0 = u_wallace_cla_csa1_csa_component_fa11_fa_and1 & u_wallace_cla_and_6_6;
  assign u_wallace_cla_csa3_csa_component_fa12_fa_xor1 = u_wallace_cla_csa3_csa_component_fa12_fa_xor0 ^ u_wallace_cla_and_5_7;
  assign u_wallace_cla_csa3_csa_component_fa12_fa_and1 = u_wallace_cla_csa3_csa_component_fa12_fa_xor0 & u_wallace_cla_and_5_7;
  assign u_wallace_cla_csa3_csa_component_fa12_fa_or0 = u_wallace_cla_csa3_csa_component_fa12_fa_and0 | u_wallace_cla_csa3_csa_component_fa12_fa_and1;
  assign u_wallace_cla_csa3_csa_component_fa13_fa_xor1 = u_wallace_cla_and_7_6 ^ u_wallace_cla_and_6_7;
  assign u_wallace_cla_csa3_csa_component_fa13_fa_and1 = u_wallace_cla_and_7_6 & u_wallace_cla_and_6_7;
  assign u_wallace_cla_csa4_csa_component_fa3_fa_xor0 = u_wallace_cla_csa2_csa_component_fa3_fa_xor1 ^ u_wallace_cla_csa2_csa_component_fa2_fa_and0;
  assign u_wallace_cla_csa4_csa_component_fa3_fa_and0 = u_wallace_cla_csa2_csa_component_fa3_fa_xor1 & u_wallace_cla_csa2_csa_component_fa2_fa_and0;
  assign u_wallace_cla_csa4_csa_component_fa4_fa_xor0 = u_wallace_cla_csa2_csa_component_fa4_fa_xor1 ^ u_wallace_cla_csa2_csa_component_fa3_fa_or0;
  assign u_wallace_cla_csa4_csa_component_fa4_fa_and0 = u_wallace_cla_csa2_csa_component_fa4_fa_xor1 & u_wallace_cla_csa2_csa_component_fa3_fa_or0;
  assign u_wallace_cla_csa4_csa_component_fa5_fa_xor0 = u_wallace_cla_csa2_csa_component_fa5_fa_xor1 ^ u_wallace_cla_csa2_csa_component_fa4_fa_or0;
  assign u_wallace_cla_csa4_csa_component_fa5_fa_and0 = u_wallace_cla_csa2_csa_component_fa5_fa_xor1 & u_wallace_cla_csa2_csa_component_fa4_fa_or0;
  assign u_wallace_cla_csa4_csa_component_fa5_fa_xor1 = u_wallace_cla_csa4_csa_component_fa5_fa_xor0 ^ u_wallace_cla_csa1_csa_component_fa4_fa_and0;
  assign u_wallace_cla_csa4_csa_component_fa5_fa_and1 = u_wallace_cla_csa4_csa_component_fa5_fa_xor0 & u_wallace_cla_csa1_csa_component_fa4_fa_and0;
  assign u_wallace_cla_csa4_csa_component_fa5_fa_or0 = u_wallace_cla_csa4_csa_component_fa5_fa_and0 | u_wallace_cla_csa4_csa_component_fa5_fa_and1;
  assign u_wallace_cla_csa4_csa_component_fa6_fa_xor0 = u_wallace_cla_csa2_csa_component_fa6_fa_xor1 ^ u_wallace_cla_csa2_csa_component_fa5_fa_or0;
  assign u_wallace_cla_csa4_csa_component_fa6_fa_and0 = u_wallace_cla_csa2_csa_component_fa6_fa_xor1 & u_wallace_cla_csa2_csa_component_fa5_fa_or0;
  assign u_wallace_cla_csa4_csa_component_fa6_fa_xor1 = u_wallace_cla_csa4_csa_component_fa6_fa_xor0 ^ u_wallace_cla_csa3_csa_component_fa6_fa_xor0;
  assign u_wallace_cla_csa4_csa_component_fa6_fa_and1 = u_wallace_cla_csa4_csa_component_fa6_fa_xor0 & u_wallace_cla_csa3_csa_component_fa6_fa_xor0;
  assign u_wallace_cla_csa4_csa_component_fa6_fa_or0 = u_wallace_cla_csa4_csa_component_fa6_fa_and0 | u_wallace_cla_csa4_csa_component_fa6_fa_and1;
  assign u_wallace_cla_csa4_csa_component_fa7_fa_xor0 = u_wallace_cla_csa2_csa_component_fa7_fa_xor1 ^ u_wallace_cla_csa2_csa_component_fa6_fa_or0;
  assign u_wallace_cla_csa4_csa_component_fa7_fa_and0 = u_wallace_cla_csa2_csa_component_fa7_fa_xor1 & u_wallace_cla_csa2_csa_component_fa6_fa_or0;
  assign u_wallace_cla_csa4_csa_component_fa7_fa_xor1 = u_wallace_cla_csa4_csa_component_fa7_fa_xor0 ^ u_wallace_cla_csa3_csa_component_fa7_fa_xor1;
  assign u_wallace_cla_csa4_csa_component_fa7_fa_and1 = u_wallace_cla_csa4_csa_component_fa7_fa_xor0 & u_wallace_cla_csa3_csa_component_fa7_fa_xor1;
  assign u_wallace_cla_csa4_csa_component_fa7_fa_or0 = u_wallace_cla_csa4_csa_component_fa7_fa_and0 | u_wallace_cla_csa4_csa_component_fa7_fa_and1;
  assign u_wallace_cla_csa4_csa_component_fa8_fa_xor0 = u_wallace_cla_csa2_csa_component_fa8_fa_xor1 ^ u_wallace_cla_csa2_csa_component_fa7_fa_or0;
  assign u_wallace_cla_csa4_csa_component_fa8_fa_and0 = u_wallace_cla_csa2_csa_component_fa8_fa_xor1 & u_wallace_cla_csa2_csa_component_fa7_fa_or0;
  assign u_wallace_cla_csa4_csa_component_fa8_fa_xor1 = u_wallace_cla_csa4_csa_component_fa8_fa_xor0 ^ u_wallace_cla_csa3_csa_component_fa8_fa_xor1;
  assign u_wallace_cla_csa4_csa_component_fa8_fa_and1 = u_wallace_cla_csa4_csa_component_fa8_fa_xor0 & u_wallace_cla_csa3_csa_component_fa8_fa_xor1;
  assign u_wallace_cla_csa4_csa_component_fa8_fa_or0 = u_wallace_cla_csa4_csa_component_fa8_fa_and0 | u_wallace_cla_csa4_csa_component_fa8_fa_and1;
  assign u_wallace_cla_csa4_csa_component_fa9_fa_xor0 = u_wallace_cla_csa2_csa_component_fa9_fa_xor1 ^ u_wallace_cla_csa2_csa_component_fa8_fa_or0;
  assign u_wallace_cla_csa4_csa_component_fa9_fa_and0 = u_wallace_cla_csa2_csa_component_fa9_fa_xor1 & u_wallace_cla_csa2_csa_component_fa8_fa_or0;
  assign u_wallace_cla_csa4_csa_component_fa9_fa_xor1 = u_wallace_cla_csa4_csa_component_fa9_fa_xor0 ^ u_wallace_cla_csa3_csa_component_fa9_fa_xor1;
  assign u_wallace_cla_csa4_csa_component_fa9_fa_and1 = u_wallace_cla_csa4_csa_component_fa9_fa_xor0 & u_wallace_cla_csa3_csa_component_fa9_fa_xor1;
  assign u_wallace_cla_csa4_csa_component_fa9_fa_or0 = u_wallace_cla_csa4_csa_component_fa9_fa_and0 | u_wallace_cla_csa4_csa_component_fa9_fa_and1;
  assign u_wallace_cla_csa4_csa_component_fa10_fa_xor0 = u_wallace_cla_csa1_csa_component_fa10_fa_xor1 ^ u_wallace_cla_csa2_csa_component_fa9_fa_or0;
  assign u_wallace_cla_csa4_csa_component_fa10_fa_and0 = u_wallace_cla_csa1_csa_component_fa10_fa_xor1 & u_wallace_cla_csa2_csa_component_fa9_fa_or0;
  assign u_wallace_cla_csa4_csa_component_fa10_fa_xor1 = u_wallace_cla_csa4_csa_component_fa10_fa_xor0 ^ u_wallace_cla_csa3_csa_component_fa10_fa_xor1;
  assign u_wallace_cla_csa4_csa_component_fa10_fa_and1 = u_wallace_cla_csa4_csa_component_fa10_fa_xor0 & u_wallace_cla_csa3_csa_component_fa10_fa_xor1;
  assign u_wallace_cla_csa4_csa_component_fa10_fa_or0 = u_wallace_cla_csa4_csa_component_fa10_fa_and0 | u_wallace_cla_csa4_csa_component_fa10_fa_and1;
  assign u_wallace_cla_csa4_csa_component_fa11_fa_xor1 = u_wallace_cla_csa1_csa_component_fa11_fa_xor1 ^ u_wallace_cla_csa3_csa_component_fa11_fa_xor1;
  assign u_wallace_cla_csa4_csa_component_fa11_fa_and1 = u_wallace_cla_csa1_csa_component_fa11_fa_xor1 & u_wallace_cla_csa3_csa_component_fa11_fa_xor1;
  assign u_wallace_cla_csa4_csa_component_fa12_fa_xor1 = u_wallace_cla_and_7_5 ^ u_wallace_cla_csa3_csa_component_fa12_fa_xor1;
  assign u_wallace_cla_csa4_csa_component_fa12_fa_and1 = u_wallace_cla_and_7_5 & u_wallace_cla_csa3_csa_component_fa12_fa_xor1;
  assign u_wallace_cla_csa5_csa_component_fa4_fa_xor0 = u_wallace_cla_csa4_csa_component_fa4_fa_xor0 ^ u_wallace_cla_csa4_csa_component_fa3_fa_and0;
  assign u_wallace_cla_csa5_csa_component_fa4_fa_and0 = u_wallace_cla_csa4_csa_component_fa4_fa_xor0 & u_wallace_cla_csa4_csa_component_fa3_fa_and0;
  assign u_wallace_cla_csa5_csa_component_fa5_fa_xor0 = u_wallace_cla_csa4_csa_component_fa5_fa_xor1 ^ u_wallace_cla_csa4_csa_component_fa4_fa_and0;
  assign u_wallace_cla_csa5_csa_component_fa5_fa_and0 = u_wallace_cla_csa4_csa_component_fa5_fa_xor1 & u_wallace_cla_csa4_csa_component_fa4_fa_and0;
  assign u_wallace_cla_csa5_csa_component_fa6_fa_xor0 = u_wallace_cla_csa4_csa_component_fa6_fa_xor1 ^ u_wallace_cla_csa4_csa_component_fa5_fa_or0;
  assign u_wallace_cla_csa5_csa_component_fa6_fa_and0 = u_wallace_cla_csa4_csa_component_fa6_fa_xor1 & u_wallace_cla_csa4_csa_component_fa5_fa_or0;
  assign u_wallace_cla_csa5_csa_component_fa7_fa_xor0 = u_wallace_cla_csa4_csa_component_fa7_fa_xor1 ^ u_wallace_cla_csa4_csa_component_fa6_fa_or0;
  assign u_wallace_cla_csa5_csa_component_fa7_fa_and0 = u_wallace_cla_csa4_csa_component_fa7_fa_xor1 & u_wallace_cla_csa4_csa_component_fa6_fa_or0;
  assign u_wallace_cla_csa5_csa_component_fa7_fa_xor1 = u_wallace_cla_csa5_csa_component_fa7_fa_xor0 ^ u_wallace_cla_csa3_csa_component_fa6_fa_and0;
  assign u_wallace_cla_csa5_csa_component_fa7_fa_and1 = u_wallace_cla_csa5_csa_component_fa7_fa_xor0 & u_wallace_cla_csa3_csa_component_fa6_fa_and0;
  assign u_wallace_cla_csa5_csa_component_fa7_fa_or0 = u_wallace_cla_csa5_csa_component_fa7_fa_and0 | u_wallace_cla_csa5_csa_component_fa7_fa_and1;
  assign u_wallace_cla_csa5_csa_component_fa8_fa_xor0 = u_wallace_cla_csa4_csa_component_fa8_fa_xor1 ^ u_wallace_cla_csa4_csa_component_fa7_fa_or0;
  assign u_wallace_cla_csa5_csa_component_fa8_fa_and0 = u_wallace_cla_csa4_csa_component_fa8_fa_xor1 & u_wallace_cla_csa4_csa_component_fa7_fa_or0;
  assign u_wallace_cla_csa5_csa_component_fa8_fa_xor1 = u_wallace_cla_csa5_csa_component_fa8_fa_xor0 ^ u_wallace_cla_csa3_csa_component_fa7_fa_or0;
  assign u_wallace_cla_csa5_csa_component_fa8_fa_and1 = u_wallace_cla_csa5_csa_component_fa8_fa_xor0 & u_wallace_cla_csa3_csa_component_fa7_fa_or0;
  assign u_wallace_cla_csa5_csa_component_fa8_fa_or0 = u_wallace_cla_csa5_csa_component_fa8_fa_and0 | u_wallace_cla_csa5_csa_component_fa8_fa_and1;
  assign u_wallace_cla_csa5_csa_component_fa9_fa_xor0 = u_wallace_cla_csa4_csa_component_fa9_fa_xor1 ^ u_wallace_cla_csa4_csa_component_fa8_fa_or0;
  assign u_wallace_cla_csa5_csa_component_fa9_fa_and0 = u_wallace_cla_csa4_csa_component_fa9_fa_xor1 & u_wallace_cla_csa4_csa_component_fa8_fa_or0;
  assign u_wallace_cla_csa5_csa_component_fa9_fa_xor1 = u_wallace_cla_csa5_csa_component_fa9_fa_xor0 ^ u_wallace_cla_csa3_csa_component_fa8_fa_or0;
  assign u_wallace_cla_csa5_csa_component_fa9_fa_and1 = u_wallace_cla_csa5_csa_component_fa9_fa_xor0 & u_wallace_cla_csa3_csa_component_fa8_fa_or0;
  assign u_wallace_cla_csa5_csa_component_fa9_fa_or0 = u_wallace_cla_csa5_csa_component_fa9_fa_and0 | u_wallace_cla_csa5_csa_component_fa9_fa_and1;
  assign u_wallace_cla_csa5_csa_component_fa10_fa_xor0 = u_wallace_cla_csa4_csa_component_fa10_fa_xor1 ^ u_wallace_cla_csa4_csa_component_fa9_fa_or0;
  assign u_wallace_cla_csa5_csa_component_fa10_fa_and0 = u_wallace_cla_csa4_csa_component_fa10_fa_xor1 & u_wallace_cla_csa4_csa_component_fa9_fa_or0;
  assign u_wallace_cla_csa5_csa_component_fa10_fa_xor1 = u_wallace_cla_csa5_csa_component_fa10_fa_xor0 ^ u_wallace_cla_csa3_csa_component_fa9_fa_or0;
  assign u_wallace_cla_csa5_csa_component_fa10_fa_and1 = u_wallace_cla_csa5_csa_component_fa10_fa_xor0 & u_wallace_cla_csa3_csa_component_fa9_fa_or0;
  assign u_wallace_cla_csa5_csa_component_fa10_fa_or0 = u_wallace_cla_csa5_csa_component_fa10_fa_and0 | u_wallace_cla_csa5_csa_component_fa10_fa_and1;
  assign u_wallace_cla_csa5_csa_component_fa11_fa_xor0 = u_wallace_cla_csa4_csa_component_fa11_fa_xor1 ^ u_wallace_cla_csa4_csa_component_fa10_fa_or0;
  assign u_wallace_cla_csa5_csa_component_fa11_fa_and0 = u_wallace_cla_csa4_csa_component_fa11_fa_xor1 & u_wallace_cla_csa4_csa_component_fa10_fa_or0;
  assign u_wallace_cla_csa5_csa_component_fa11_fa_xor1 = u_wallace_cla_csa5_csa_component_fa11_fa_xor0 ^ u_wallace_cla_csa3_csa_component_fa10_fa_or0;
  assign u_wallace_cla_csa5_csa_component_fa11_fa_and1 = u_wallace_cla_csa5_csa_component_fa11_fa_xor0 & u_wallace_cla_csa3_csa_component_fa10_fa_or0;
  assign u_wallace_cla_csa5_csa_component_fa11_fa_or0 = u_wallace_cla_csa5_csa_component_fa11_fa_and0 | u_wallace_cla_csa5_csa_component_fa11_fa_and1;
  assign u_wallace_cla_csa5_csa_component_fa12_fa_xor0 = u_wallace_cla_csa4_csa_component_fa12_fa_xor1 ^ u_wallace_cla_csa4_csa_component_fa11_fa_and1;
  assign u_wallace_cla_csa5_csa_component_fa12_fa_and0 = u_wallace_cla_csa4_csa_component_fa12_fa_xor1 & u_wallace_cla_csa4_csa_component_fa11_fa_and1;
  assign u_wallace_cla_csa5_csa_component_fa12_fa_xor1 = u_wallace_cla_csa5_csa_component_fa12_fa_xor0 ^ u_wallace_cla_csa3_csa_component_fa11_fa_or0;
  assign u_wallace_cla_csa5_csa_component_fa12_fa_and1 = u_wallace_cla_csa5_csa_component_fa12_fa_xor0 & u_wallace_cla_csa3_csa_component_fa11_fa_or0;
  assign u_wallace_cla_csa5_csa_component_fa12_fa_or0 = u_wallace_cla_csa5_csa_component_fa12_fa_and0 | u_wallace_cla_csa5_csa_component_fa12_fa_and1;
  assign u_wallace_cla_csa5_csa_component_fa13_fa_xor0 = u_wallace_cla_csa3_csa_component_fa13_fa_xor1 ^ u_wallace_cla_csa4_csa_component_fa12_fa_and1;
  assign u_wallace_cla_csa5_csa_component_fa13_fa_and0 = u_wallace_cla_csa3_csa_component_fa13_fa_xor1 & u_wallace_cla_csa4_csa_component_fa12_fa_and1;
  assign u_wallace_cla_csa5_csa_component_fa13_fa_xor1 = u_wallace_cla_csa5_csa_component_fa13_fa_xor0 ^ u_wallace_cla_csa3_csa_component_fa12_fa_or0;
  assign u_wallace_cla_csa5_csa_component_fa13_fa_and1 = u_wallace_cla_csa5_csa_component_fa13_fa_xor0 & u_wallace_cla_csa3_csa_component_fa12_fa_or0;
  assign u_wallace_cla_csa5_csa_component_fa13_fa_or0 = u_wallace_cla_csa5_csa_component_fa13_fa_and0 | u_wallace_cla_csa5_csa_component_fa13_fa_and1;
  assign u_wallace_cla_csa5_csa_component_fa14_fa_xor1 = u_wallace_cla_and_7_7 ^ u_wallace_cla_csa3_csa_component_fa13_fa_and1;
  assign u_wallace_cla_csa5_csa_component_fa14_fa_and1 = u_wallace_cla_and_7_7 & u_wallace_cla_csa3_csa_component_fa13_fa_and1;
  assign u_wallace_cla_u_cla16_and0_2_0_1_0 = u_wallace_cla_csa2_csa_component_fa2_fa_xor0 & u_wallace_cla_and_0_0;
  assign u_wallace_cla_u_cla16_and0_3_0_1_1 = u_wallace_cla_csa4_csa_component_fa3_fa_xor0 & u_wallace_cla_csa0_csa_component_fa1_fa_xor0;
  assign u_wallace_cla_u_cla16_and0_3_1_1_2 = u_wallace_cla_csa4_csa_component_fa3_fa_xor0 & u_wallace_cla_csa0_csa_component_fa1_fa_xor0;
  assign u_wallace_cla_u_cla16_pg_logic5_pg_logic_or0 = u_wallace_cla_csa5_csa_component_fa5_fa_xor0 | u_wallace_cla_csa5_csa_component_fa4_fa_and0;
  assign u_wallace_cla_u_cla16_pg_logic5_pg_logic_and0 = u_wallace_cla_csa5_csa_component_fa5_fa_xor0 & u_wallace_cla_csa5_csa_component_fa4_fa_and0;
  assign u_wallace_cla_u_cla16_pg_logic5_pg_logic_xor0 = u_wallace_cla_csa5_csa_component_fa5_fa_xor0 ^ u_wallace_cla_csa5_csa_component_fa4_fa_and0;
  assign u_wallace_cla_u_cla16_pg_logic6_pg_logic_or0 = u_wallace_cla_csa5_csa_component_fa6_fa_xor0 | u_wallace_cla_csa5_csa_component_fa5_fa_and0;
  assign u_wallace_cla_u_cla16_pg_logic6_pg_logic_and0 = u_wallace_cla_csa5_csa_component_fa6_fa_xor0 & u_wallace_cla_csa5_csa_component_fa5_fa_and0;
  assign u_wallace_cla_u_cla16_pg_logic6_pg_logic_xor0 = u_wallace_cla_csa5_csa_component_fa6_fa_xor0 ^ u_wallace_cla_csa5_csa_component_fa5_fa_and0;
  assign u_wallace_cla_u_cla16_xor6 = u_wallace_cla_u_cla16_pg_logic6_pg_logic_xor0 ^ u_wallace_cla_u_cla16_pg_logic5_pg_logic_and0;
  assign u_wallace_cla_u_cla16_and1_2_0_1_3 = u_wallace_cla_u_cla16_pg_logic6_pg_logic_or0 & u_wallace_cla_csa5_csa_component_fa4_fa_xor0;
  assign u_wallace_cla_u_cla16_and1_2_2_0_4 = u_wallace_cla_u_cla16_pg_logic5_pg_logic_and0 & u_wallace_cla_u_cla16_pg_logic6_pg_logic_or0;
  assign u_wallace_cla_u_cla16_or1_2_2_0 = u_wallace_cla_u_cla16_pg_logic6_pg_logic_and0 | u_wallace_cla_u_cla16_and1_2_2_0_4;
  assign u_wallace_cla_u_cla16_pg_logic7_pg_logic_or0 = u_wallace_cla_csa5_csa_component_fa7_fa_xor1 | u_wallace_cla_csa5_csa_component_fa6_fa_and0;
  assign u_wallace_cla_u_cla16_pg_logic7_pg_logic_and0 = u_wallace_cla_csa5_csa_component_fa7_fa_xor1 & u_wallace_cla_csa5_csa_component_fa6_fa_and0;
  assign u_wallace_cla_u_cla16_pg_logic7_pg_logic_xor0 = u_wallace_cla_csa5_csa_component_fa7_fa_xor1 ^ u_wallace_cla_csa5_csa_component_fa6_fa_and0;
  assign u_wallace_cla_u_cla16_xor7 = u_wallace_cla_u_cla16_pg_logic7_pg_logic_xor0 ^ u_wallace_cla_u_cla16_or1_2_2_0;
  assign u_wallace_cla_u_cla16_and1_3_0_1_5 = u_wallace_cla_u_cla16_pg_logic7_pg_logic_or0 & u_wallace_cla_u_cla16_pg_logic5_pg_logic_or0;
  assign u_wallace_cla_u_cla16_and1_3_1_1_6 = u_wallace_cla_u_cla16_pg_logic7_pg_logic_or0 & u_wallace_cla_u_cla16_pg_logic5_pg_logic_or0;
  assign u_wallace_cla_u_cla16_and1_3_2_0_7 = u_wallace_cla_u_cla16_pg_logic5_pg_logic_and0 & u_wallace_cla_u_cla16_pg_logic7_pg_logic_or0;
  assign u_wallace_cla_u_cla16_and1_3_2_1_8 = u_wallace_cla_u_cla16_and1_3_2_0_7 & u_wallace_cla_u_cla16_pg_logic6_pg_logic_or0;
  assign u_wallace_cla_u_cla16_and1_3_3_0_9 = u_wallace_cla_u_cla16_pg_logic6_pg_logic_and0 & u_wallace_cla_u_cla16_pg_logic7_pg_logic_or0;
  assign u_wallace_cla_u_cla16_orred1_3_3__2_1 = u_wallace_cla_u_cla16_and1_3_2_1_8 | u_wallace_cla_u_cla16_and1_3_3_0_9;
  assign u_wallace_cla_u_cla16_or1_3_3_2 = u_wallace_cla_u_cla16_pg_logic7_pg_logic_and0 | u_wallace_cla_u_cla16_orred1_3_3__2_1;
  assign u_wallace_cla_u_cla16_pg_logic8_pg_logic_or0 = u_wallace_cla_csa5_csa_component_fa8_fa_xor1 | u_wallace_cla_csa5_csa_component_fa7_fa_or0;
  assign u_wallace_cla_u_cla16_pg_logic8_pg_logic_and0 = u_wallace_cla_csa5_csa_component_fa8_fa_xor1 & u_wallace_cla_csa5_csa_component_fa7_fa_or0;
  assign u_wallace_cla_u_cla16_pg_logic8_pg_logic_xor0 = u_wallace_cla_csa5_csa_component_fa8_fa_xor1 ^ u_wallace_cla_csa5_csa_component_fa7_fa_or0;
  assign u_wallace_cla_u_cla16_xor8 = u_wallace_cla_u_cla16_pg_logic8_pg_logic_xor0 ^ u_wallace_cla_u_cla16_or1_3_3_2;
  assign u_wallace_cla_u_cla16_and2_0_0_0_10 = u_wallace_cla_u_cla16_or1_3_3_2 & u_wallace_cla_u_cla16_pg_logic8_pg_logic_or0;
  assign u_wallace_cla_u_cla16_or2_0_0_3 = u_wallace_cla_u_cla16_pg_logic8_pg_logic_and0 | u_wallace_cla_u_cla16_and2_0_0_0_10;
  assign u_wallace_cla_u_cla16_pg_logic9_pg_logic_or0 = u_wallace_cla_csa5_csa_component_fa9_fa_xor1 | u_wallace_cla_csa5_csa_component_fa8_fa_or0;
  assign u_wallace_cla_u_cla16_pg_logic9_pg_logic_and0 = u_wallace_cla_csa5_csa_component_fa9_fa_xor1 & u_wallace_cla_csa5_csa_component_fa8_fa_or0;
  assign u_wallace_cla_u_cla16_pg_logic9_pg_logic_xor0 = u_wallace_cla_csa5_csa_component_fa9_fa_xor1 ^ u_wallace_cla_csa5_csa_component_fa8_fa_or0;
  assign u_wallace_cla_u_cla16_xor9 = u_wallace_cla_u_cla16_pg_logic9_pg_logic_xor0 ^ u_wallace_cla_u_cla16_or2_0_0_3;
  assign u_wallace_cla_u_cla16_and2_1_0_0_11 = u_wallace_cla_u_cla16_or1_3_3_2 & u_wallace_cla_u_cla16_pg_logic9_pg_logic_or0;
  assign u_wallace_cla_u_cla16_and2_1_0_1_12 = u_wallace_cla_u_cla16_and2_1_0_0_11 & u_wallace_cla_u_cla16_pg_logic8_pg_logic_or0;
  assign u_wallace_cla_u_cla16_and2_1_1_0_13 = u_wallace_cla_u_cla16_pg_logic8_pg_logic_and0 & u_wallace_cla_u_cla16_pg_logic9_pg_logic_or0;
  assign u_wallace_cla_u_cla16_orred2_1_1__0_4 = u_wallace_cla_u_cla16_and2_1_0_1_12 | u_wallace_cla_u_cla16_and2_1_1_0_13;
  assign u_wallace_cla_u_cla16_or2_1_1_5 = u_wallace_cla_u_cla16_pg_logic9_pg_logic_and0 | u_wallace_cla_u_cla16_orred2_1_1__0_4;
  assign u_wallace_cla_u_cla16_pg_logic10_pg_logic_or0 = u_wallace_cla_csa5_csa_component_fa10_fa_xor1 | u_wallace_cla_csa5_csa_component_fa9_fa_or0;
  assign u_wallace_cla_u_cla16_pg_logic10_pg_logic_and0 = u_wallace_cla_csa5_csa_component_fa10_fa_xor1 & u_wallace_cla_csa5_csa_component_fa9_fa_or0;
  assign u_wallace_cla_u_cla16_pg_logic10_pg_logic_xor0 = u_wallace_cla_csa5_csa_component_fa10_fa_xor1 ^ u_wallace_cla_csa5_csa_component_fa9_fa_or0;
  assign u_wallace_cla_u_cla16_xor10 = u_wallace_cla_u_cla16_pg_logic10_pg_logic_xor0 ^ u_wallace_cla_u_cla16_or2_1_1_5;
  assign u_wallace_cla_u_cla16_and2_2_0_0_14 = u_wallace_cla_u_cla16_or1_3_3_2 & u_wallace_cla_u_cla16_pg_logic9_pg_logic_or0;
  assign u_wallace_cla_u_cla16_and2_2_0_1_15 = u_wallace_cla_u_cla16_pg_logic10_pg_logic_or0 & u_wallace_cla_u_cla16_pg_logic8_pg_logic_or0;
  assign u_wallace_cla_u_cla16_and2_2_0_2_16 = u_wallace_cla_u_cla16_and2_2_0_0_14 & u_wallace_cla_u_cla16_and2_2_0_1_15;
  assign u_wallace_cla_u_cla16_and2_2_1_0_17 = u_wallace_cla_u_cla16_pg_logic8_pg_logic_and0 & u_wallace_cla_u_cla16_pg_logic10_pg_logic_or0;
  assign u_wallace_cla_u_cla16_and2_2_1_1_18 = u_wallace_cla_u_cla16_and2_2_1_0_17 & u_wallace_cla_u_cla16_pg_logic9_pg_logic_or0;
  assign u_wallace_cla_u_cla16_and2_2_2_0_19 = u_wallace_cla_u_cla16_pg_logic9_pg_logic_and0 & u_wallace_cla_u_cla16_pg_logic10_pg_logic_or0;
  assign u_wallace_cla_u_cla16_orred2_2_2__0_6 = u_wallace_cla_u_cla16_and2_2_0_2_16 | u_wallace_cla_u_cla16_and2_2_1_1_18;
  assign u_wallace_cla_u_cla16_orred2_2_2__1_7 = u_wallace_cla_u_cla16_orred2_2_2__0_6 | u_wallace_cla_u_cla16_and2_2_2_0_19;
  assign u_wallace_cla_u_cla16_or2_2_2_8 = u_wallace_cla_u_cla16_pg_logic10_pg_logic_and0 | u_wallace_cla_u_cla16_orred2_2_2__1_7;
  assign u_wallace_cla_u_cla16_pg_logic11_pg_logic_or0 = u_wallace_cla_csa5_csa_component_fa11_fa_xor1 | u_wallace_cla_csa5_csa_component_fa10_fa_or0;
  assign u_wallace_cla_u_cla16_pg_logic11_pg_logic_and0 = u_wallace_cla_csa5_csa_component_fa11_fa_xor1 & u_wallace_cla_csa5_csa_component_fa10_fa_or0;
  assign u_wallace_cla_u_cla16_pg_logic11_pg_logic_xor0 = u_wallace_cla_csa5_csa_component_fa11_fa_xor1 ^ u_wallace_cla_csa5_csa_component_fa10_fa_or0;
  assign u_wallace_cla_u_cla16_xor11 = u_wallace_cla_u_cla16_pg_logic11_pg_logic_xor0 ^ u_wallace_cla_u_cla16_or2_2_2_8;
  assign u_wallace_cla_u_cla16_and2_3_0_0_20 = u_wallace_cla_u_cla16_or1_3_3_2 & u_wallace_cla_u_cla16_pg_logic10_pg_logic_or0;
  assign u_wallace_cla_u_cla16_and2_3_0_1_21 = u_wallace_cla_u_cla16_pg_logic11_pg_logic_or0 & u_wallace_cla_u_cla16_pg_logic9_pg_logic_or0;
  assign u_wallace_cla_u_cla16_and2_3_0_2_22 = u_wallace_cla_u_cla16_and2_3_0_0_20 & u_wallace_cla_u_cla16_and2_3_0_1_21;
  assign u_wallace_cla_u_cla16_and2_3_0_3_23 = u_wallace_cla_u_cla16_and2_3_0_2_22 & u_wallace_cla_u_cla16_pg_logic8_pg_logic_or0;
  assign u_wallace_cla_u_cla16_and2_3_1_0_24 = u_wallace_cla_u_cla16_pg_logic8_pg_logic_and0 & u_wallace_cla_u_cla16_pg_logic10_pg_logic_or0;
  assign u_wallace_cla_u_cla16_and2_3_1_1_25 = u_wallace_cla_u_cla16_pg_logic11_pg_logic_or0 & u_wallace_cla_u_cla16_pg_logic9_pg_logic_or0;
  assign u_wallace_cla_u_cla16_and2_3_1_2_26 = u_wallace_cla_u_cla16_and2_3_1_0_24 & u_wallace_cla_u_cla16_and2_3_1_1_25;
  assign u_wallace_cla_u_cla16_and2_3_2_0_27 = u_wallace_cla_u_cla16_pg_logic9_pg_logic_and0 & u_wallace_cla_u_cla16_pg_logic11_pg_logic_or0;
  assign u_wallace_cla_u_cla16_and2_3_2_1_28 = u_wallace_cla_u_cla16_and2_3_2_0_27 & u_wallace_cla_u_cla16_pg_logic10_pg_logic_or0;
  assign u_wallace_cla_u_cla16_and2_3_3_0_29 = u_wallace_cla_u_cla16_pg_logic10_pg_logic_and0 & u_wallace_cla_u_cla16_pg_logic11_pg_logic_or0;
  assign u_wallace_cla_u_cla16_orred2_3_3__0_9 = u_wallace_cla_u_cla16_and2_3_0_3_23 | u_wallace_cla_u_cla16_and2_3_2_1_28;
  assign u_wallace_cla_u_cla16_orred2_3_3__1_10 = u_wallace_cla_u_cla16_and2_3_1_2_26 | u_wallace_cla_u_cla16_and2_3_3_0_29;
  assign u_wallace_cla_u_cla16_orred2_3_3__2_11 = u_wallace_cla_u_cla16_orred2_3_3__0_9 | u_wallace_cla_u_cla16_orred2_3_3__1_10;
  assign u_wallace_cla_u_cla16_or2_3_3_12 = u_wallace_cla_u_cla16_pg_logic11_pg_logic_and0 | u_wallace_cla_u_cla16_orred2_3_3__2_11;
  assign u_wallace_cla_u_cla16_pg_logic12_pg_logic_or0 = u_wallace_cla_csa5_csa_component_fa12_fa_xor1 | u_wallace_cla_csa5_csa_component_fa11_fa_or0;
  assign u_wallace_cla_u_cla16_pg_logic12_pg_logic_and0 = u_wallace_cla_csa5_csa_component_fa12_fa_xor1 & u_wallace_cla_csa5_csa_component_fa11_fa_or0;
  assign u_wallace_cla_u_cla16_pg_logic12_pg_logic_xor0 = u_wallace_cla_csa5_csa_component_fa12_fa_xor1 ^ u_wallace_cla_csa5_csa_component_fa11_fa_or0;
  assign u_wallace_cla_u_cla16_xor12 = u_wallace_cla_u_cla16_pg_logic12_pg_logic_xor0 ^ u_wallace_cla_u_cla16_or2_3_3_12;
  assign u_wallace_cla_u_cla16_and3_0_0_0_30 = u_wallace_cla_u_cla16_or2_3_3_12 & u_wallace_cla_u_cla16_pg_logic12_pg_logic_or0;
  assign u_wallace_cla_u_cla16_or3_0_0_13 = u_wallace_cla_u_cla16_pg_logic12_pg_logic_and0 | u_wallace_cla_u_cla16_and3_0_0_0_30;
  assign u_wallace_cla_u_cla16_pg_logic13_pg_logic_or0 = u_wallace_cla_csa5_csa_component_fa13_fa_xor1 | u_wallace_cla_csa5_csa_component_fa12_fa_or0;
  assign u_wallace_cla_u_cla16_pg_logic13_pg_logic_and0 = u_wallace_cla_csa5_csa_component_fa13_fa_xor1 & u_wallace_cla_csa5_csa_component_fa12_fa_or0;
  assign u_wallace_cla_u_cla16_pg_logic13_pg_logic_xor0 = u_wallace_cla_csa5_csa_component_fa13_fa_xor1 ^ u_wallace_cla_csa5_csa_component_fa12_fa_or0;
  assign u_wallace_cla_u_cla16_xor13 = u_wallace_cla_u_cla16_pg_logic13_pg_logic_xor0 ^ u_wallace_cla_u_cla16_or3_0_0_13;
  assign u_wallace_cla_u_cla16_and3_1_0_0_31 = u_wallace_cla_u_cla16_or2_3_3_12 & u_wallace_cla_u_cla16_pg_logic13_pg_logic_or0;
  assign u_wallace_cla_u_cla16_and3_1_0_1_32 = u_wallace_cla_u_cla16_and3_1_0_0_31 & u_wallace_cla_u_cla16_pg_logic12_pg_logic_or0;
  assign u_wallace_cla_u_cla16_and3_1_1_0_33 = u_wallace_cla_u_cla16_pg_logic12_pg_logic_and0 & u_wallace_cla_u_cla16_pg_logic13_pg_logic_or0;
  assign u_wallace_cla_u_cla16_orred3_1_1__0_14 = u_wallace_cla_u_cla16_and3_1_0_1_32 | u_wallace_cla_u_cla16_and3_1_1_0_33;
  assign u_wallace_cla_u_cla16_or3_1_1_15 = u_wallace_cla_u_cla16_pg_logic13_pg_logic_and0 | u_wallace_cla_u_cla16_orred3_1_1__0_14;
  assign u_wallace_cla_u_cla16_pg_logic14_pg_logic_or0 = u_wallace_cla_csa5_csa_component_fa14_fa_xor1 | u_wallace_cla_csa5_csa_component_fa13_fa_or0;
  assign u_wallace_cla_u_cla16_pg_logic14_pg_logic_and0 = u_wallace_cla_csa5_csa_component_fa14_fa_xor1 & u_wallace_cla_csa5_csa_component_fa13_fa_or0;
  assign u_wallace_cla_u_cla16_pg_logic14_pg_logic_xor0 = u_wallace_cla_csa5_csa_component_fa14_fa_xor1 ^ u_wallace_cla_csa5_csa_component_fa13_fa_or0;
  assign u_wallace_cla_u_cla16_xor14 = u_wallace_cla_u_cla16_pg_logic14_pg_logic_xor0 ^ u_wallace_cla_u_cla16_or3_1_1_15;
  assign u_wallace_cla_u_cla16_and3_2_0_0_34 = u_wallace_cla_u_cla16_or2_3_3_12 & u_wallace_cla_u_cla16_pg_logic13_pg_logic_or0;
  assign u_wallace_cla_u_cla16_and3_2_0_1_35 = u_wallace_cla_u_cla16_pg_logic14_pg_logic_or0 & u_wallace_cla_u_cla16_pg_logic12_pg_logic_or0;
  assign u_wallace_cla_u_cla16_and3_2_0_2_36 = u_wallace_cla_u_cla16_and3_2_0_0_34 & u_wallace_cla_u_cla16_and3_2_0_1_35;
  assign u_wallace_cla_u_cla16_and3_2_1_0_37 = u_wallace_cla_u_cla16_pg_logic12_pg_logic_and0 & u_wallace_cla_u_cla16_pg_logic14_pg_logic_or0;
  assign u_wallace_cla_u_cla16_and3_2_1_1_38 = u_wallace_cla_u_cla16_and3_2_1_0_37 & u_wallace_cla_u_cla16_pg_logic13_pg_logic_or0;
  assign u_wallace_cla_u_cla16_and3_2_2_0_39 = u_wallace_cla_u_cla16_pg_logic13_pg_logic_and0 & u_wallace_cla_u_cla16_pg_logic14_pg_logic_or0;
  assign u_wallace_cla_u_cla16_orred3_2_2__0_16 = u_wallace_cla_u_cla16_and3_2_0_2_36 | u_wallace_cla_u_cla16_and3_2_1_1_38;
  assign u_wallace_cla_u_cla16_orred3_2_2__1_17 = u_wallace_cla_u_cla16_orred3_2_2__0_16 | u_wallace_cla_u_cla16_and3_2_2_0_39;
  assign u_wallace_cla_u_cla16_or3_2_2_18 = u_wallace_cla_u_cla16_pg_logic14_pg_logic_and0 | u_wallace_cla_u_cla16_orred3_2_2__1_17;
  assign u_wallace_cla_u_cla16_xor15 = u_wallace_cla_csa5_csa_component_fa14_fa_and1 ^ u_wallace_cla_u_cla16_or3_2_2_18;
  assign u_wallace_cla_u_cla16_and3_3_0_0_40 = u_wallace_cla_u_cla16_or2_3_3_12 & u_wallace_cla_u_cla16_pg_logic14_pg_logic_or0;
  assign u_wallace_cla_u_cla16_and3_3_0_1_41 = u_wallace_cla_csa5_csa_component_fa14_fa_and1 & u_wallace_cla_u_cla16_pg_logic13_pg_logic_or0;
  assign u_wallace_cla_u_cla16_and3_3_0_2_42 = u_wallace_cla_u_cla16_and3_3_0_0_40 & u_wallace_cla_u_cla16_and3_3_0_1_41;
  assign u_wallace_cla_u_cla16_and3_3_0_3_43 = u_wallace_cla_u_cla16_and3_3_0_2_42 & u_wallace_cla_u_cla16_pg_logic12_pg_logic_or0;
  assign u_wallace_cla_u_cla16_and3_3_1_0_44 = u_wallace_cla_u_cla16_pg_logic12_pg_logic_and0 & u_wallace_cla_u_cla16_pg_logic14_pg_logic_or0;
  assign u_wallace_cla_u_cla16_and3_3_1_1_45 = u_wallace_cla_csa5_csa_component_fa14_fa_and1 & u_wallace_cla_u_cla16_pg_logic13_pg_logic_or0;
  assign u_wallace_cla_u_cla16_and3_3_1_2_46 = u_wallace_cla_u_cla16_and3_3_1_0_44 & u_wallace_cla_u_cla16_and3_3_1_1_45;
  assign u_wallace_cla_u_cla16_and3_3_2_0_47 = u_wallace_cla_u_cla16_pg_logic13_pg_logic_and0 & u_wallace_cla_csa5_csa_component_fa14_fa_and1;
  assign u_wallace_cla_u_cla16_and3_3_2_1_48 = u_wallace_cla_u_cla16_and3_3_2_0_47 & u_wallace_cla_u_cla16_pg_logic14_pg_logic_or0;
  assign u_wallace_cla_u_cla16_and3_3_3_0_49 = u_wallace_cla_u_cla16_pg_logic14_pg_logic_and0 & u_wallace_cla_csa5_csa_component_fa14_fa_and1;
  assign u_wallace_cla_u_cla16_orred3_3_3__0_19 = u_wallace_cla_u_cla16_and3_3_0_3_43 | u_wallace_cla_u_cla16_and3_3_2_1_48;
  assign u_wallace_cla_u_cla16_orred3_3_3__1_20 = u_wallace_cla_u_cla16_and3_3_1_2_46 | u_wallace_cla_u_cla16_and3_3_3_0_49;
  assign u_wallace_cla_u_cla16_orred3_3_3__2_21 = u_wallace_cla_u_cla16_orred3_3_3__0_19 | u_wallace_cla_u_cla16_orred3_3_3__1_20;

  assign u_wallace_cla_out[0] = u_wallace_cla_and_0_0;
  assign u_wallace_cla_out[1] = u_wallace_cla_csa0_csa_component_fa1_fa_xor0;
  assign u_wallace_cla_out[2] = u_wallace_cla_csa2_csa_component_fa2_fa_xor0;
  assign u_wallace_cla_out[3] = u_wallace_cla_csa4_csa_component_fa3_fa_xor0;
  assign u_wallace_cla_out[4] = u_wallace_cla_csa5_csa_component_fa4_fa_xor0;
  assign u_wallace_cla_out[5] = u_wallace_cla_u_cla16_pg_logic5_pg_logic_xor0;
  assign u_wallace_cla_out[6] = u_wallace_cla_u_cla16_xor6;
  assign u_wallace_cla_out[7] = u_wallace_cla_u_cla16_xor7;
  assign u_wallace_cla_out[8] = u_wallace_cla_u_cla16_xor8;
  assign u_wallace_cla_out[9] = u_wallace_cla_u_cla16_xor9;
  assign u_wallace_cla_out[10] = u_wallace_cla_u_cla16_xor10;
  assign u_wallace_cla_out[11] = u_wallace_cla_u_cla16_xor11;
  assign u_wallace_cla_out[12] = u_wallace_cla_u_cla16_xor12;
  assign u_wallace_cla_out[13] = u_wallace_cla_u_cla16_xor13;
  assign u_wallace_cla_out[14] = u_wallace_cla_u_cla16_xor14;
  assign u_wallace_cla_out[15] = u_wallace_cla_u_cla16_xor15;
endmodule